magic
tech sky130A
magscale 1 2
timestamp 1761874473
<< nwell >>
rect -1309 1035 -550 1356
rect -4130 -191 -3351 130
rect -2302 -195 -1513 126
rect -1108 -193 -269 128
rect 812 -193 1533 128
rect -4178 -1715 -3245 -1394
rect -2184 -1709 -1427 -1388
rect -994 -1711 -243 -1390
rect 774 -1713 1573 -1392
rect -1373 -2895 -550 -2574
<< pwell >>
rect -1209 795 -487 977
rect -4153 -431 -3451 -249
rect -2345 -431 -1681 -249
rect -1133 -433 -369 -251
rect 775 -433 1433 -251
rect -4137 -1955 -3345 -1773
rect -2295 -1949 -1494 -1767
rect -963 -1951 -343 -1769
rect 791 -1953 1473 -1771
rect -1273 -3135 -507 -2953
<< viali >>
rect -2344 989 -2300 1033
rect -1770 989 -1674 1085
rect -1327 989 -1287 1029
rect -3307 -237 -3263 -193
rect -2906 -237 -2810 -141
rect -2554 -237 -2514 -197
rect -1442 -241 -1392 -191
rect -1049 -254 -985 -190
rect -347 -239 -313 -205
rect 532 -237 566 -203
rect 871 -233 905 -199
rect 1396 -233 1430 -199
rect 2108 -281 2159 -229
rect -3372 -1761 -3328 -1717
rect -2800 -1761 -2704 -1665
rect -2444 -1761 -2404 -1721
rect -1188 -1755 -1138 -1705
rect -963 -1770 -899 -1706
rect -321 -1751 -287 -1717
rect 490 -1757 524 -1723
rect 883 -1759 917 -1725
rect 1436 -1759 1470 -1725
rect 2148 -1779 2199 -1727
rect -2319 -2941 -2275 -2897
rect -1834 -2941 -1738 -2845
rect -1478 -2941 -1438 -2901
<< metal1 >>
rect -4656 1335 -2467 1366
rect -1057 1335 -507 1366
rect -4653 140 -4622 1335
rect -1770 1091 -1674 1136
rect -1776 1085 -1668 1091
rect -2350 1033 -2294 1039
rect -2882 989 -2344 1033
rect -2300 989 -2244 1033
rect -2350 983 -2294 989
rect -1776 983 -1770 1085
rect -1674 983 -1668 1085
rect -1520 983 -1514 1035
rect -1462 1029 -1456 1035
rect -1333 1029 -1281 1035
rect -1462 989 -1327 1029
rect -1287 989 -1192 1029
rect -1462 983 -1456 989
rect -1333 983 -1281 989
rect -1770 902 -1674 908
rect -1059 785 -545 816
rect -4363 716 -4357 768
rect -4305 757 -4299 768
rect -4305 726 -2462 757
rect -4305 716 -4299 726
rect -4656 109 -3603 140
rect -4379 -110 -4348 109
rect -2221 105 -1765 136
rect -1015 107 -518 138
rect 865 107 1281 138
rect -4396 -162 -4390 -110
rect -4338 -162 -4332 -110
rect -2912 -141 -2804 -135
rect -3258 -187 -3206 -183
rect -3313 -189 -3206 -187
rect -3313 -193 -3258 -189
rect -3370 -237 -3307 -193
rect -3263 -237 -3258 -193
rect -3313 -241 -3258 -237
rect -2990 -237 -2906 -141
rect -2810 -237 -2712 -141
rect -1448 -190 -1386 -185
rect -1055 -190 -979 -184
rect -1448 -191 -1442 -190
rect -1390 -191 -1384 -190
rect -2564 -197 -2558 -191
rect -2506 -197 -2500 -191
rect -2626 -237 -2558 -197
rect -2506 -237 -2448 -197
rect -3313 -243 -3206 -241
rect -2912 -243 -2804 -237
rect -2564 -243 -2558 -237
rect -2506 -243 -2500 -237
rect -1525 -241 -1442 -191
rect -1390 -241 -1349 -191
rect -1448 -242 -1442 -241
rect -1390 -242 -1384 -241
rect -3258 -247 -3206 -243
rect -1448 -247 -1386 -242
rect -1072 -254 -1049 -190
rect -985 -205 -504 -190
rect 522 -194 574 -188
rect -353 -205 -307 -199
rect 865 -199 911 -187
rect 1390 -199 1436 -193
rect -985 -239 -347 -205
rect -313 -239 -213 -205
rect 463 -237 522 -203
rect 574 -237 631 -203
rect 865 -233 871 -199
rect 905 -233 1396 -199
rect 1430 -233 1471 -199
rect 2102 -229 2165 -217
rect -985 -254 -504 -239
rect -353 -245 -307 -239
rect 865 -245 911 -233
rect 522 -252 574 -246
rect -1055 -260 -979 -254
rect 1081 -262 1115 -233
rect 1390 -239 1436 -233
rect 1072 -268 1124 -262
rect 2071 -280 2108 -229
rect 2102 -281 2108 -280
rect 2159 -280 2559 -229
rect 2159 -281 2165 -280
rect 2102 -293 2165 -281
rect 1072 -326 1124 -320
rect -4099 -435 -3583 -404
rect -2197 -439 -1757 -408
rect -1019 -437 -521 -406
rect 867 -437 1284 -406
rect -4665 -458 -4613 -452
rect -4613 -500 -4129 -469
rect -4665 -516 -4613 -510
rect -4391 -984 -4339 -978
rect -4391 -1042 -4339 -1036
rect -4381 -1384 -4350 -1042
rect -4381 -1415 -3497 -1384
rect -2180 -1407 -1676 -1378
rect -4381 -1797 -4350 -1415
rect -2180 -1444 -2151 -1407
rect -917 -1411 -495 -1380
rect 915 -1411 1329 -1380
rect -672 -1506 -620 -1500
rect -672 -1564 -620 -1558
rect 1096 -1548 1148 -1542
rect -2806 -1665 -2698 -1659
rect -3776 -1717 -3716 -1712
rect -3378 -1717 -3322 -1711
rect -3776 -1718 -3372 -1717
rect -3716 -1761 -3372 -1718
rect -3328 -1761 -3204 -1717
rect -2870 -1761 -2800 -1665
rect -2704 -1761 -2636 -1665
rect -1194 -1704 -1132 -1699
rect -1196 -1705 -1190 -1704
rect -1138 -1705 -1132 -1704
rect -2422 -1715 -2370 -1709
rect -2450 -1721 -2422 -1715
rect -2514 -1761 -2444 -1721
rect -2370 -1761 -2330 -1721
rect -1281 -1755 -1190 -1705
rect -1138 -1755 -1077 -1705
rect -969 -1706 -893 -1700
rect -1196 -1756 -1190 -1755
rect -1138 -1756 -1132 -1755
rect -1194 -1761 -1132 -1756
rect -3716 -1778 -3204 -1761
rect -2806 -1767 -2698 -1761
rect -2450 -1767 -2422 -1761
rect -2422 -1773 -2370 -1767
rect -986 -1770 -963 -1706
rect -899 -1714 -752 -1706
rect -899 -1766 -840 -1714
rect -788 -1766 -752 -1714
rect -663 -1717 -629 -1564
rect 1096 -1606 1148 -1600
rect -327 -1717 -281 -1711
rect -663 -1751 -321 -1717
rect -287 -1751 -237 -1717
rect 476 -1723 482 -1714
rect 534 -1723 540 -1714
rect -327 -1757 -281 -1751
rect 441 -1757 482 -1723
rect 534 -1757 571 -1723
rect 871 -1725 929 -1719
rect 1105 -1725 1139 -1606
rect 1430 -1725 1476 -1719
rect 2148 -1721 2199 -1681
rect 476 -1766 482 -1757
rect 534 -1766 540 -1757
rect 871 -1759 883 -1725
rect 917 -1759 1436 -1725
rect 1470 -1759 1519 -1725
rect 2142 -1727 2205 -1721
rect 871 -1765 929 -1759
rect -899 -1770 -752 -1766
rect -969 -1776 -893 -1770
rect -840 -1772 -788 -1770
rect -3776 -1784 -3716 -1778
rect 1105 -1794 1139 -1759
rect 1430 -1765 1476 -1759
rect 2107 -1778 2148 -1727
rect 2142 -1779 2148 -1778
rect 2199 -1728 2241 -1727
rect 2199 -1779 2575 -1728
rect 2142 -1785 2205 -1779
rect -4391 -1803 -4339 -1797
rect -4391 -1861 -4339 -1855
rect 1096 -1800 1148 -1794
rect 2148 -1819 2199 -1785
rect 1096 -1858 1148 -1852
rect -4095 -1959 -3494 -1928
rect -2109 -1953 -1679 -1922
rect -945 -1955 -495 -1924
rect 909 -1957 1321 -1926
rect -4561 -1982 -4509 -1976
rect -4509 -2024 -4113 -1993
rect -4561 -2040 -4509 -2034
rect -3336 -2219 -3284 -2213
rect -3336 -2277 -3284 -2271
rect -3325 -2564 -3294 -2277
rect -3325 -2595 -2506 -2564
rect -1139 -2597 -565 -2566
rect -1840 -2845 -1732 -2839
rect -2325 -2897 -2269 -2891
rect -2820 -2941 -2319 -2897
rect -2275 -2941 -2200 -2897
rect -1890 -2941 -1834 -2845
rect -1736 -2941 -1670 -2845
rect -2325 -2947 -2269 -2941
rect -1840 -2947 -1732 -2941
rect -1628 -2947 -1622 -2895
rect -1570 -2901 -1564 -2895
rect -1484 -2901 -1432 -2895
rect -1570 -2941 -1478 -2901
rect -1438 -2941 -1366 -2901
rect -1570 -2947 -1564 -2941
rect -1484 -2947 -1432 -2941
rect -1124 -3139 -567 -3108
rect -3633 -3214 -3627 -3162
rect -3575 -3173 -3569 -3162
rect -3575 -3204 -2398 -3173
rect -3575 -3214 -3569 -3204
<< via1 >>
rect -1770 989 -1674 1004
rect -1770 908 -1674 989
rect -1514 983 -1462 1035
rect -4357 716 -4305 768
rect -4390 -162 -4338 -110
rect -3258 -241 -3206 -189
rect -2906 -237 -2810 -141
rect -1442 -191 -1390 -190
rect -2558 -197 -2506 -191
rect -2558 -237 -2554 -197
rect -2554 -237 -2514 -197
rect -2514 -237 -2506 -197
rect -2558 -243 -2506 -237
rect -1442 -241 -1392 -191
rect -1392 -241 -1390 -191
rect -1442 -242 -1390 -241
rect 522 -203 574 -194
rect 522 -237 532 -203
rect 532 -237 566 -203
rect 566 -237 574 -203
rect 522 -246 574 -237
rect 1072 -320 1124 -268
rect -4665 -510 -4613 -458
rect -4391 -1036 -4339 -984
rect -672 -1558 -620 -1506
rect -3776 -1778 -3716 -1718
rect -2800 -1761 -2704 -1665
rect -1190 -1705 -1138 -1704
rect -2422 -1721 -2370 -1715
rect -2422 -1761 -2404 -1721
rect -2404 -1761 -2370 -1721
rect -1190 -1755 -1188 -1705
rect -1188 -1755 -1138 -1705
rect -1190 -1756 -1138 -1755
rect -2422 -1767 -2370 -1761
rect -840 -1766 -788 -1714
rect 1096 -1600 1148 -1548
rect 482 -1723 534 -1714
rect 482 -1757 490 -1723
rect 490 -1757 524 -1723
rect 524 -1757 534 -1723
rect 482 -1766 534 -1757
rect -4391 -1855 -4339 -1803
rect 1096 -1852 1148 -1800
rect -4561 -2034 -4509 -1982
rect -3336 -2271 -3284 -2219
rect -1832 -2941 -1738 -2845
rect -1738 -2941 -1736 -2845
rect -1622 -2947 -1570 -2895
rect -3627 -3214 -3575 -3162
<< metal2 >>
rect -1514 1035 -1462 1041
rect -1774 1004 -1514 1029
rect -1776 908 -1770 1004
rect -1674 989 -1514 1004
rect -1674 908 -1668 989
rect -1514 977 -1462 983
rect -4357 768 -4305 774
rect -4971 727 -4357 758
rect -4971 -1992 -4940 727
rect -4357 710 -4305 716
rect -1770 534 -1674 908
rect -2906 438 -1386 534
rect -4390 -110 -4338 -104
rect -4390 -168 -4338 -162
rect -2906 -141 -2810 438
rect -4671 -510 -4665 -458
rect -4613 -510 -4607 -458
rect -4654 -1992 -4623 -510
rect -4380 -984 -4349 -168
rect -3264 -241 -3258 -189
rect -3206 -241 -3200 -189
rect -3254 -522 -3210 -241
rect -4397 -1036 -4391 -984
rect -4339 -1036 -4333 -984
rect -3289 -998 -3174 -522
rect -2906 -740 -2810 -237
rect -2558 -191 -2506 -185
rect -2558 -249 -2506 -243
rect -2552 -613 -2512 -249
rect -2396 -613 -2340 -606
rect -2552 -615 -2338 -613
rect -2552 -671 -2396 -615
rect -2340 -671 -2338 -615
rect -2552 -673 -2338 -671
rect -2396 -680 -2340 -673
rect -2906 -836 -2345 -740
rect -3289 -1094 -2704 -998
rect -3289 -1097 -3174 -1094
rect -2800 -1665 -2704 -1094
rect -3774 -1718 -3718 -1711
rect -3782 -1778 -3776 -1718
rect -3716 -1778 -3710 -1718
rect -3774 -1785 -3718 -1778
rect -4397 -1855 -4391 -1803
rect -4339 -1855 -4333 -1803
rect -4567 -1992 -4561 -1982
rect -4973 -2023 -4561 -1992
rect -4971 -2451 -4940 -2023
rect -4654 -2025 -4623 -2023
rect -4567 -2034 -4561 -2023
rect -4509 -2034 -4503 -1982
rect -4380 -2230 -4349 -1855
rect -3342 -2230 -3336 -2219
rect -4380 -2261 -3336 -2230
rect -3342 -2271 -3336 -2261
rect -3284 -2271 -3278 -2219
rect -2800 -2286 -2704 -1761
rect -2446 -1715 -2345 -836
rect -2072 -744 -1976 438
rect -1441 -184 -1391 438
rect -1442 -190 -1390 -184
rect -1442 -248 -1390 -242
rect 516 -246 522 -194
rect 574 -246 580 -194
rect -2072 -840 -1136 -744
rect -1040 -840 -1031 -744
rect 531 -1211 565 -246
rect 1066 -320 1072 -268
rect 1124 -320 1130 -268
rect 747 -613 807 -604
rect 1081 -626 1115 -320
rect 807 -661 1116 -626
rect 747 -682 807 -673
rect 1081 -847 1115 -661
rect 1068 -856 1128 -847
rect 1068 -925 1128 -916
rect -2446 -1767 -2422 -1715
rect -2370 -1767 -2345 -1715
rect -2446 -1791 -2345 -1767
rect -1928 -1312 -1302 -1216
rect -1206 -1312 -1190 -1216
rect 382 -1246 438 -1239
rect 531 -1245 1139 -1211
rect -664 -1248 440 -1246
rect -664 -1304 382 -1248
rect 438 -1304 440 -1248
rect -664 -1306 440 -1304
rect -1928 -2286 -1832 -1312
rect -663 -1506 -629 -1306
rect 382 -1313 438 -1306
rect -678 -1558 -672 -1506
rect -620 -1558 -614 -1506
rect 1105 -1548 1139 -1245
rect 1090 -1600 1096 -1548
rect 1148 -1600 1154 -1548
rect -1190 -1704 -1138 -1698
rect 482 -1714 534 -1708
rect -1190 -1762 -1138 -1756
rect -1189 -2286 -1139 -1762
rect -846 -1766 -840 -1714
rect -788 -1723 -782 -1714
rect -788 -1757 482 -1723
rect -788 -1766 -782 -1757
rect 482 -1772 534 -1766
rect 1090 -1852 1096 -1800
rect 1148 -1852 1154 -1800
rect -719 -2224 -710 -2164
rect -650 -2177 -641 -2164
rect 1105 -2177 1139 -1852
rect -650 -2211 1139 -2177
rect -650 -2224 -641 -2211
rect -2800 -2382 -1138 -2286
rect -4971 -2482 -4245 -2451
rect -4971 -2488 -4940 -2482
rect -4276 -3172 -4245 -2482
rect -1832 -2845 -1736 -2382
rect -1622 -2895 -1570 -2889
rect -1736 -2941 -1622 -2901
rect -1832 -2947 -1736 -2941
rect -1622 -2953 -1570 -2947
rect -3627 -3162 -3575 -3156
rect -4276 -3203 -3627 -3172
rect -3627 -3220 -3575 -3214
<< via2 >>
rect -2396 -671 -2340 -615
rect -3774 -1776 -3718 -1720
rect -1136 -840 -1040 -744
rect 747 -673 807 -613
rect 1068 -916 1128 -856
rect -1302 -1312 -1206 -1216
rect 382 -1304 438 -1248
rect -710 -2224 -650 -2164
<< metal3 >>
rect -2401 -613 -2335 -610
rect 742 -613 812 -608
rect -2401 -615 747 -613
rect -2401 -671 -2396 -615
rect -2340 -671 747 -615
rect -2401 -673 747 -671
rect 807 -673 910 -613
rect -2401 -676 -2335 -673
rect 742 -678 812 -673
rect -1141 -744 -1035 -739
rect -1141 -840 -1136 -744
rect -1040 -840 -1035 -744
rect -1141 -845 -1035 -840
rect -1136 -964 -1040 -845
rect 1063 -856 1133 -851
rect 1063 -916 1068 -856
rect 1128 -916 1133 -856
rect 1063 -921 1133 -916
rect -1307 -1216 -1201 -1211
rect -1136 -1216 -1040 -1116
rect -1307 -1312 -1302 -1216
rect -1206 -1312 -1040 -1216
rect 377 -1246 443 -1243
rect 1068 -1246 1128 -921
rect 377 -1248 1128 -1246
rect 377 -1304 382 -1248
rect 438 -1304 1128 -1248
rect 377 -1306 1128 -1304
rect 377 -1309 443 -1306
rect -1307 -1317 -1201 -1312
rect -1134 -1314 -1042 -1312
rect -3779 -1720 -3713 -1715
rect -3779 -1776 -3774 -1720
rect -3718 -1776 -3713 -1720
rect -3779 -1781 -3713 -1776
rect -3776 -2164 -3716 -1781
rect -715 -2164 -645 -2159
rect -3776 -2224 -710 -2164
rect -650 -2224 -645 -2164
rect -715 -2229 -645 -2224
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_3 ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1760154773
transform 1 0 -4144 0 1 -1976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_5
timestamp 1760154773
transform 1 0 -596 0 1 -3158
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_6
timestamp 1760154773
transform 1 0 -4160 0 1 -452
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_8
timestamp 1760154773
transform 1 0 -576 0 1 768
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_8  x1 ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 -2498 0 1 774
box -38 -48 1510 592
use sky130_fd_sc_hd__nand2_8  x2
timestamp 1704896540
transform 1 0 -3634 0 1 -452
box -38 -48 1510 592
use sky130_fd_sc_hd__nand2_8  x3
timestamp 1704896540
transform 1 0 -3528 0 1 -1976
box -38 -48 1510 592
use sky130_fd_sc_hd__nand2_8  x4
timestamp 1704896540
transform 1 0 -2562 0 1 -3156
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_8  x5 ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 -1796 0 1 -456
box -38 -48 866 592
use sky130_fd_sc_hd__inv_8  x6
timestamp 1704896540
transform 1 0 -1710 0 1 -1970
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_8  x7 ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 -552 0 1 -454
box -38 -48 1510 592
use sky130_fd_sc_hd__nor2_8  x8
timestamp 1704896540
transform 1 0 -526 0 1 -1972
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_8  x9 ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 1290 0 1 -1974
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  x10
timestamp 1704896540
transform 1 0 1250 0 1 -454
box -38 -48 1142 592
<< labels >>
rlabel space -4656 1335 -507 1366 7 VPWR
port 2 w
rlabel metal2 -4971 727 -4357 758 7 VGND
port 3 w
rlabel metal1 -2820 -2941 -2319 -2897 7 ENABLE
port 1 w
rlabel metal1 2159 -280 2559 -229 3 Qn
port 5 e
rlabel metal3 -1136 -1312 -1040 -1116 1 C1
port 7 n
rlabel metal3 -1136 -964 -1040 -840 5 C2
port 8 s
rlabel metal1 -2882 989 -2838 1033 7 ENABLE
port 1 w
rlabel metal1 2199 -1779 2575 -1728 3 Q
port 4 e
<< end >>
