magic
tech sky130A
magscale 1 2
timestamp 1761264907
<< pwell >>
rect 19573 21763 19797 21849
rect 19573 21637 19659 21763
rect 19573 21551 20249 21637
rect 20163 21417 20249 21551
<< metal1 >>
rect 22688 29512 22694 29572
rect 22754 29512 22760 29572
rect 22694 27323 22754 29512
rect 25694 27982 25746 27988
rect 25694 27924 25746 27930
rect 22527 27272 25403 27323
rect 17180 27264 17232 27270
rect 17180 27206 17232 27212
rect 17184 24789 17228 27206
rect 17184 24745 17780 24789
rect 25352 23542 25403 27272
rect 24992 23491 25403 23542
rect 8303 22919 8309 23090
rect 8480 23055 11110 23090
rect 8480 23033 13987 23055
rect 8480 22975 16615 23033
rect 8480 22953 13987 22975
rect 8480 22919 11110 22953
rect 25697 21957 25743 27924
rect 25053 21911 25743 21957
rect 19567 21434 20013 21465
rect 17140 20811 17146 20863
rect 17198 20859 17204 20863
rect 17198 20815 17518 20859
rect 17198 20811 17204 20815
<< via1 >>
rect 22694 29512 22754 29572
rect 25694 27930 25746 27982
rect 17180 27212 17232 27264
rect 8309 22919 8480 23090
rect 17146 20811 17198 20863
<< metal2 >>
rect 23246 35964 23306 35966
rect 23239 35908 23248 35964
rect 23304 35908 23313 35964
rect 22694 35838 22754 35840
rect 22687 35782 22696 35838
rect 22752 35782 22761 35838
rect 17176 30308 17236 30317
rect 17176 30239 17236 30248
rect 17184 27264 17228 30239
rect 22694 29572 22754 35782
rect 22694 29506 22754 29512
rect 23246 27979 23306 35908
rect 25688 27979 25694 27982
rect 22947 27933 25694 27979
rect 25688 27930 25694 27933
rect 25746 27930 25752 27982
rect 17174 27212 17180 27264
rect 17232 27212 17238 27264
rect 8309 23090 8480 23096
rect 2668 22919 2677 23090
rect 2848 22919 8309 23090
rect 8309 22913 8480 22919
rect 10382 22483 10391 22641
rect 10549 22618 13185 22641
rect 10549 22595 14070 22618
rect 10549 22578 15117 22595
rect 10549 22546 16822 22578
rect 10549 22529 15117 22546
rect 10549 22506 14070 22529
rect 10549 22483 13185 22506
rect 16027 20807 16036 20867
rect 16096 20859 16105 20867
rect 17146 20863 17198 20869
rect 16096 20815 17146 20859
rect 16096 20807 16105 20815
rect 17146 20805 17198 20811
<< via2 >>
rect 23248 35908 23304 35964
rect 22696 35782 22752 35838
rect 17176 30248 17236 30308
rect 2677 22919 2848 23090
rect 10391 22483 10549 22641
rect 16036 20807 16096 20867
<< metal3 >>
rect 22686 39578 22692 39642
rect 22756 39578 22762 39642
rect 23238 39578 23244 39642
rect 23308 39578 23314 39642
rect 22694 35843 22754 39578
rect 23246 35969 23306 39578
rect 23243 35964 23309 35969
rect 23243 35908 23248 35964
rect 23304 35908 23309 35964
rect 23243 35903 23309 35908
rect 22691 35838 22757 35843
rect 22691 35782 22696 35838
rect 22752 35782 22757 35838
rect 22691 35777 22757 35782
rect 17174 31994 17238 32000
rect 17174 31924 17238 31930
rect 17176 30313 17236 31924
rect 17171 30308 17241 30313
rect 17171 30248 17176 30308
rect 17236 30248 17241 30308
rect 17171 30243 17241 30248
rect 16034 27620 16098 27626
rect 16034 27550 16098 27556
rect 226 23090 480 23226
rect 2672 23090 2853 23095
rect 226 22919 279 23090
rect 450 22919 2677 23090
rect 2848 22919 2853 23090
rect 226 22800 480 22919
rect 2672 22914 2853 22919
rect 10386 22641 10554 22646
rect 2683 22483 2689 22641
rect 2847 22483 10391 22641
rect 10549 22483 10554 22641
rect 10386 22478 10554 22483
rect 16036 20872 16096 27550
rect 20726 23256 20732 23258
rect 20078 23196 20732 23256
rect 20726 23194 20732 23196
rect 20796 23194 20802 23258
rect 19479 22921 20067 22991
rect 16031 20867 16101 20872
rect 16031 20807 16036 20867
rect 16096 20807 16101 20867
rect 16031 20802 16101 20807
rect 18779 19871 18849 19877
rect 19479 19871 19549 22921
rect 19997 22854 20067 22921
rect 18849 19801 19549 19871
rect 18779 19795 18849 19801
<< via3 >>
rect 22692 39578 22756 39642
rect 23244 39578 23308 39642
rect 17174 31930 17238 31994
rect 16034 27556 16098 27620
rect 279 22919 450 23090
rect 2689 22483 2847 22641
rect 20732 23194 20796 23258
rect 18779 19801 18849 19871
<< metal4 >>
rect 6134 44952 6194 45152
rect 6686 44952 6746 45152
rect 7238 44952 7298 45152
rect 7790 44952 7850 45152
rect 8342 44952 8402 45152
rect 8894 44952 8954 45152
rect 9446 44952 9506 45152
rect 9998 44952 10058 45152
rect 10550 44952 10610 45152
rect 11102 44952 11162 45152
rect 11654 44952 11714 45152
rect 12206 44952 12266 45152
rect 12758 44952 12818 45152
rect 13310 44952 13370 45152
rect 13862 44952 13922 45152
rect 14414 44952 14474 45152
rect 14966 44952 15026 45152
rect 15518 44952 15578 45152
rect 16070 44952 16130 45152
rect 16622 44952 16682 45152
rect 17174 44952 17234 45152
rect 17726 44952 17786 45152
rect 18278 44952 18338 45152
rect 18830 44952 18890 45152
rect 19382 44952 19442 45152
rect 19934 44952 19994 45152
rect 20486 44952 20546 45152
rect 21038 44952 21098 45152
rect 200 23090 600 44152
rect 200 22919 279 23090
rect 450 22919 600 23090
rect 200 1000 600 22919
rect 800 22641 1200 44152
rect 19945 44119 20698 44122
rect 17233 44100 20698 44119
rect 21590 44100 21650 45152
rect 17233 44040 21650 44100
rect 17233 44021 20698 44040
rect 21590 44034 21650 44040
rect 17233 34731 17331 44021
rect 19945 44019 20698 44021
rect 15695 34633 17331 34731
rect 18627 43124 20773 43151
rect 18627 43104 21332 43124
rect 22142 43104 22202 45152
rect 18627 43044 22202 43104
rect 18627 43025 21332 43044
rect 18627 42997 20773 43025
rect 16036 27621 16096 34633
rect 18627 33727 18781 42997
rect 22694 39643 22754 45152
rect 23246 39643 23306 45152
rect 23798 44952 23858 45152
rect 24350 44952 24410 45152
rect 24902 44952 24962 45152
rect 25454 44952 25514 45152
rect 26006 44952 26066 45152
rect 26558 44952 26618 45152
rect 27110 44952 27170 45152
rect 27662 44952 27722 45152
rect 28214 44952 28274 45152
rect 28766 44952 28826 45152
rect 29318 44952 29378 45152
rect 22691 39642 22757 39643
rect 22691 39578 22692 39642
rect 22756 39578 22757 39642
rect 22691 39577 22757 39578
rect 23243 39642 23309 39643
rect 23243 39578 23244 39642
rect 23308 39578 23309 39642
rect 23243 39577 23309 39578
rect 16755 33573 18781 33727
rect 17176 31995 17236 33573
rect 17173 31994 17239 31995
rect 17173 31930 17174 31994
rect 17238 31930 17239 31994
rect 17173 31929 17239 31930
rect 16033 27620 16099 27621
rect 16033 27556 16034 27620
rect 16098 27556 16099 27620
rect 16033 27555 16099 27556
rect 20731 23258 20797 23259
rect 20731 23194 20732 23258
rect 20796 23194 20797 23258
rect 20731 23193 20797 23194
rect 2688 22641 2848 22642
rect 800 22483 2689 22641
rect 2847 22483 2848 22641
rect 800 1000 1200 22483
rect 2688 22482 2848 22483
rect 18778 19871 18850 19872
rect 18778 19801 18779 19871
rect 18849 19801 18850 19871
rect 18778 19800 18850 19801
rect 20734 19830 20794 23193
rect 18779 18690 18849 19800
rect 20734 19770 21068 19830
rect 21008 19080 21068 19770
rect 18694 10638 18874 18690
rect 20902 14014 21082 19080
rect 20902 13834 30542 14014
rect 18694 10458 26678 10638
rect 3314 0 3494 200
rect 7178 0 7358 200
rect 11042 0 11222 200
rect 14906 0 15086 200
rect 18770 0 18950 200
rect 22634 0 22814 200
rect 26498 0 26678 10458
rect 30362 0 30542 13834
use layout_mod  layout_mod_0 ~/Downloads
timestamp 1761264109
transform 1 0 20372 0 1 23756
box -3936 -3276 4733 2024
<< labels >>
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 29318 44952 29378 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 28214 44952 28274 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 30362 0 30542 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26498 0 26678 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22634 0 22814 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18770 0 18950 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 14906 0 15086 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 11042 0 11222 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 7178 0 7358 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 3314 0 3494 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 27662 44952 27722 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 27110 44952 27170 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 26006 44952 26066 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 25454 44952 25514 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 24902 44952 24962 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 23798 44952 23858 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23246 44952 23306 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22694 44952 22754 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21590 44952 21650 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 21038 44952 21098 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 20486 44952 20546 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 19382 44952 19442 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 9998 44952 10058 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 9446 44952 9506 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 8342 44952 8402 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 7790 44952 7850 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 7238 44952 7298 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 6134 44952 6194 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 14414 44952 14474 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 13862 44952 13922 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 12758 44952 12818 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 12206 44952 12266 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 11654 44952 11714 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 10550 44952 10610 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 18830 44952 18890 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 18278 44952 18338 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 17174 44952 17234 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 16622 44952 16682 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 16070 44952 16130 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 14966 44952 15026 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 600 44152 1 FreeSans 400 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 800 1000 1200 44152 1 FreeSans 400 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
