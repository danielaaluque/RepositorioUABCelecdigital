magic
tech sky130A
magscale 1 2
timestamp 1762480118
<< metal1 >>
rect 27656 23396 27662 23456
rect 27722 23396 27728 23456
rect 27662 21650 27722 23396
rect 15333 21649 27722 21650
rect 15283 21590 27722 21649
rect 15283 20916 15333 21590
rect 23246 21122 23306 21128
rect 22688 21034 22694 21094
rect 22754 21093 22813 21094
rect 22754 21034 22859 21093
rect 18074 20634 18254 20640
rect 17382 20454 18074 20634
rect 18074 20448 18254 20454
rect 15298 20352 15304 20448
rect 15400 20352 15636 20448
rect 22813 19654 22859 21034
rect 22633 19608 22859 19654
rect 23036 21062 23246 21122
rect 23036 18256 23076 21062
rect 23246 21056 23306 21062
rect 22630 18216 23076 18256
rect 11742 18042 12142 18048
rect 12142 17642 14546 18042
rect 11742 17636 12142 17642
rect 15411 17400 15821 17494
rect 18002 17492 18182 17498
rect 17444 17312 18002 17492
rect 18002 17306 18182 17312
rect 15327 17115 15333 17167
rect 15385 17162 15391 17167
rect 15385 17119 15478 17162
rect 15385 17115 15391 17119
<< via1 >>
rect 27662 23396 27722 23456
rect 22694 21034 22754 21094
rect 18074 20454 18254 20634
rect 15304 20352 15400 20448
rect 23246 21062 23306 21122
rect 11742 17642 12142 18042
rect 18002 17312 18182 17492
rect 15333 17115 15385 17167
<< metal2 >>
rect 27662 28252 27722 28254
rect 27655 28196 27664 28252
rect 27720 28196 27729 28252
rect 27110 27624 27170 27626
rect 27103 27568 27112 27624
rect 27168 27568 27177 27624
rect 27110 23558 27170 27568
rect 14620 23498 27170 23558
rect 9005 18042 9395 18046
rect 9000 18037 11742 18042
rect 9000 17647 9005 18037
rect 9395 17647 11742 18037
rect 9000 17642 11742 17647
rect 12142 17642 12148 18042
rect 9005 17638 9395 17642
rect 14621 17163 14664 23498
rect 27662 23456 27722 28196
rect 27662 23390 27722 23396
rect 23246 22780 23306 22782
rect 22694 22772 22754 22774
rect 22687 22716 22696 22772
rect 22752 22716 22761 22772
rect 23239 22724 23248 22780
rect 23304 22724 23313 22780
rect 22694 21094 22754 22716
rect 23246 21122 23306 22724
rect 23240 21062 23246 21122
rect 23306 21062 23312 21122
rect 22694 21028 22754 21034
rect 19919 20634 20089 20638
rect 18068 20454 18074 20634
rect 18254 20629 20094 20634
rect 18254 20459 19919 20629
rect 20089 20459 20094 20629
rect 18254 20454 20094 20459
rect 15304 20448 15400 20454
rect 19919 20450 20089 20454
rect 14777 20352 14786 20448
rect 14882 20352 15304 20448
rect 15304 20346 15400 20352
rect 17996 17312 18002 17492
rect 18182 17487 19426 17492
rect 18182 17317 19251 17487
rect 19421 17317 19430 17487
rect 18182 17312 19426 17317
rect 15333 17167 15385 17173
rect 14621 17120 15333 17163
rect 15333 17109 15385 17115
<< via2 >>
rect 27664 28196 27720 28252
rect 27112 27568 27168 27624
rect 9005 17647 9395 18037
rect 22696 22716 22752 22772
rect 23248 22724 23304 22780
rect 19919 20459 20089 20629
rect 14786 20352 14882 20448
rect 19251 17317 19421 17487
<< metal3 >>
rect 6126 44440 6132 44504
rect 6196 44440 6202 44504
rect 17724 44468 17788 44474
rect 2094 43664 2100 43728
rect 2164 43726 2170 43728
rect 6134 43726 6194 44440
rect 17172 44438 17236 44444
rect 6678 44290 6684 44354
rect 6748 44290 6754 44354
rect 6686 43726 6746 44290
rect 7230 44276 7236 44340
rect 7300 44276 7306 44340
rect 7782 44290 7788 44354
rect 7852 44290 7858 44354
rect 8340 44342 8404 44348
rect 7238 43726 7298 44276
rect 7790 43726 7850 44290
rect 8340 44272 8404 44278
rect 8886 44276 8892 44340
rect 8956 44276 8962 44340
rect 8342 43726 8402 44272
rect 8894 43726 8954 44276
rect 9438 44244 9444 44308
rect 9508 44244 9514 44308
rect 9990 44290 9996 44354
rect 10060 44290 10066 44354
rect 10542 44302 10548 44366
rect 10612 44302 10618 44366
rect 9446 43726 9506 44244
rect 9998 43726 10058 44290
rect 10550 43726 10610 44302
rect 11094 44276 11100 44340
rect 11164 44276 11170 44340
rect 11102 43726 11162 44276
rect 11646 44250 11652 44314
rect 11716 44250 11722 44314
rect 12198 44278 12204 44342
rect 12268 44278 12274 44342
rect 11654 43726 11714 44250
rect 12206 43726 12266 44278
rect 12750 44262 12756 44326
rect 12820 44262 12826 44326
rect 13302 44290 13308 44354
rect 13372 44290 13378 44354
rect 13854 44308 13860 44372
rect 13924 44308 13930 44372
rect 12758 43726 12818 44262
rect 13310 43726 13370 44290
rect 13862 43726 13922 44308
rect 14406 44290 14412 44354
rect 14476 44290 14482 44354
rect 14414 43726 14474 44290
rect 14958 44260 14964 44324
rect 15028 44260 15034 44324
rect 15510 44302 15516 44366
rect 15580 44302 15586 44366
rect 16062 44330 16068 44394
rect 16132 44330 16138 44394
rect 16614 44364 16620 44428
rect 16684 44364 16690 44428
rect 17724 44398 17788 44404
rect 18270 44400 18276 44464
rect 18340 44400 18346 44464
rect 17172 44368 17236 44374
rect 14966 43726 15026 44260
rect 15518 43726 15578 44302
rect 16070 43726 16130 44330
rect 16622 43726 16682 44364
rect 17174 43726 17234 44368
rect 17726 43726 17786 44398
rect 2164 43666 17786 43726
rect 2164 43664 2170 43666
rect 18278 41618 18338 44400
rect 18822 44384 18828 44448
rect 18892 44384 18898 44448
rect 18830 42212 18890 44384
rect 27660 44168 27724 44174
rect 27102 44102 27108 44166
rect 27172 44102 27178 44166
rect 18830 42152 23306 42212
rect 18278 41558 22754 41618
rect 22694 22777 22754 41558
rect 23246 22785 23306 42152
rect 27110 27629 27170 44102
rect 27660 44098 27724 44104
rect 27662 28257 27722 44098
rect 27659 28252 27725 28257
rect 27659 28196 27664 28252
rect 27720 28196 27725 28252
rect 27659 28191 27725 28196
rect 27107 27624 27173 27629
rect 27107 27568 27112 27624
rect 27168 27568 27173 27624
rect 27107 27563 27173 27568
rect 23243 22780 23309 22785
rect 22691 22772 22757 22777
rect 22691 22716 22696 22772
rect 22752 22716 22757 22772
rect 23243 22724 23248 22780
rect 23304 22724 23309 22780
rect 23243 22719 23309 22724
rect 22691 22711 22757 22716
rect 19914 20629 30542 20634
rect 19914 20459 19919 20629
rect 20089 20459 30542 20629
rect 19914 20454 30542 20459
rect 14781 20448 14887 20453
rect 13870 20352 14786 20448
rect 14882 20352 14887 20448
rect 200 20124 6221 20142
rect 200 19758 220 20124
rect 574 20086 6221 20124
rect 13877 20086 14159 20352
rect 14781 20347 14887 20352
rect 574 19804 14159 20086
rect 574 19758 6221 19804
rect 200 19748 6221 19758
rect 200 19742 600 19748
rect 3099 18042 3497 18047
rect 3098 18041 9400 18042
rect 3098 17643 3099 18041
rect 3497 18037 9400 18041
rect 3497 17647 9005 18037
rect 9395 17647 9400 18037
rect 3497 17643 9400 17647
rect 3098 17642 9400 17643
rect 3099 17637 3497 17642
rect 19246 17487 26678 17492
rect 19246 17317 19251 17487
rect 19421 17317 26678 17487
rect 19246 17312 26678 17317
rect 26498 1059 26678 17312
rect 26493 881 26499 1059
rect 26677 881 26683 1059
rect 30362 921 30542 20454
rect 26498 880 26678 881
rect 30357 743 30363 921
rect 30541 743 30547 921
rect 30362 742 30542 743
<< via3 >>
rect 6132 44440 6196 44504
rect 2100 43664 2164 43728
rect 6684 44290 6748 44354
rect 7236 44276 7300 44340
rect 7788 44290 7852 44354
rect 8340 44278 8404 44342
rect 8892 44276 8956 44340
rect 9444 44244 9508 44308
rect 9996 44290 10060 44354
rect 10548 44302 10612 44366
rect 11100 44276 11164 44340
rect 11652 44250 11716 44314
rect 12204 44278 12268 44342
rect 12756 44262 12820 44326
rect 13308 44290 13372 44354
rect 13860 44308 13924 44372
rect 14412 44290 14476 44354
rect 14964 44260 15028 44324
rect 15516 44302 15580 44366
rect 16068 44330 16132 44394
rect 16620 44364 16684 44428
rect 17172 44374 17236 44438
rect 17724 44404 17788 44468
rect 18276 44400 18340 44464
rect 18828 44384 18892 44448
rect 27108 44102 27172 44166
rect 27660 44104 27724 44168
rect 220 19758 574 20124
rect 3099 17643 3497 18041
rect 26499 881 26677 1059
rect 30363 743 30541 921
<< metal4 >>
rect 6134 44505 6194 45152
rect 6131 44504 6197 44505
rect 6131 44440 6132 44504
rect 6196 44440 6197 44504
rect 6131 44439 6197 44440
rect 6686 44355 6746 45152
rect 6683 44354 6749 44355
rect 6683 44290 6684 44354
rect 6748 44290 6749 44354
rect 7238 44341 7298 45152
rect 7790 44355 7850 45152
rect 7787 44354 7853 44355
rect 6683 44289 6749 44290
rect 7235 44340 7301 44341
rect 7235 44276 7236 44340
rect 7300 44276 7301 44340
rect 7787 44290 7788 44354
rect 7852 44290 7853 44354
rect 8342 44343 8402 45152
rect 7787 44289 7853 44290
rect 8339 44342 8405 44343
rect 8339 44278 8340 44342
rect 8404 44278 8405 44342
rect 8894 44341 8954 45152
rect 8339 44277 8405 44278
rect 8891 44340 8957 44341
rect 7235 44275 7301 44276
rect 8891 44276 8892 44340
rect 8956 44276 8957 44340
rect 9446 44309 9506 45152
rect 9998 44355 10058 45152
rect 10550 44367 10610 45152
rect 10547 44366 10613 44367
rect 9995 44354 10061 44355
rect 8891 44275 8957 44276
rect 9443 44308 9509 44309
rect 9443 44244 9444 44308
rect 9508 44244 9509 44308
rect 9995 44290 9996 44354
rect 10060 44290 10061 44354
rect 10547 44302 10548 44366
rect 10612 44302 10613 44366
rect 11102 44341 11162 45152
rect 10547 44301 10613 44302
rect 11099 44340 11165 44341
rect 9995 44289 10061 44290
rect 11099 44276 11100 44340
rect 11164 44276 11165 44340
rect 11654 44315 11714 45152
rect 12206 44343 12266 45152
rect 12203 44342 12269 44343
rect 11099 44275 11165 44276
rect 11651 44314 11717 44315
rect 11651 44250 11652 44314
rect 11716 44250 11717 44314
rect 12203 44278 12204 44342
rect 12268 44278 12269 44342
rect 12758 44327 12818 45152
rect 13310 44355 13370 45152
rect 13862 44373 13922 45152
rect 13859 44372 13925 44373
rect 13307 44354 13373 44355
rect 12203 44277 12269 44278
rect 12755 44326 12821 44327
rect 12755 44262 12756 44326
rect 12820 44262 12821 44326
rect 13307 44290 13308 44354
rect 13372 44290 13373 44354
rect 13859 44308 13860 44372
rect 13924 44308 13925 44372
rect 14414 44355 14474 45152
rect 13859 44307 13925 44308
rect 14411 44354 14477 44355
rect 13307 44289 13373 44290
rect 14411 44290 14412 44354
rect 14476 44290 14477 44354
rect 14966 44325 15026 45152
rect 15518 44367 15578 45152
rect 16070 44395 16130 45152
rect 16622 44429 16682 45152
rect 17174 44439 17234 45152
rect 17726 44469 17786 45152
rect 17723 44468 17789 44469
rect 17171 44438 17237 44439
rect 16619 44428 16685 44429
rect 16067 44394 16133 44395
rect 15515 44366 15581 44367
rect 14411 44289 14477 44290
rect 14963 44324 15029 44325
rect 12755 44261 12821 44262
rect 14963 44260 14964 44324
rect 15028 44260 15029 44324
rect 15515 44302 15516 44366
rect 15580 44302 15581 44366
rect 16067 44330 16068 44394
rect 16132 44330 16133 44394
rect 16619 44364 16620 44428
rect 16684 44364 16685 44428
rect 17171 44374 17172 44438
rect 17236 44374 17237 44438
rect 17723 44404 17724 44468
rect 17788 44404 17789 44468
rect 18278 44465 18338 45152
rect 17723 44403 17789 44404
rect 18275 44464 18341 44465
rect 18275 44400 18276 44464
rect 18340 44400 18341 44464
rect 18830 44449 18890 45152
rect 19382 44952 19442 45152
rect 19934 44952 19994 45152
rect 20486 44952 20546 45152
rect 21038 44952 21098 45152
rect 21590 44952 21650 45152
rect 22142 44952 22202 45152
rect 22694 44952 22754 45152
rect 23246 44952 23306 45152
rect 23798 44952 23858 45152
rect 24350 44952 24410 45152
rect 24902 44952 24962 45152
rect 25454 44952 25514 45152
rect 26006 44952 26066 45152
rect 26558 44952 26618 45152
rect 18275 44399 18341 44400
rect 18827 44448 18893 44449
rect 18827 44384 18828 44448
rect 18892 44384 18893 44448
rect 18827 44383 18893 44384
rect 17171 44373 17237 44374
rect 16619 44363 16685 44364
rect 16067 44329 16133 44330
rect 15515 44301 15581 44302
rect 14963 44259 15029 44260
rect 11651 44249 11717 44250
rect 9443 44243 9509 44244
rect 27110 44167 27170 45152
rect 27662 44169 27722 45152
rect 28214 44952 28274 45152
rect 28766 44952 28826 45152
rect 29318 44952 29378 45152
rect 27659 44168 27725 44169
rect 27107 44166 27173 44167
rect 200 20124 600 44152
rect 200 19758 220 20124
rect 574 19758 600 20124
rect 200 1000 600 19758
rect 800 43726 1200 44152
rect 27107 44102 27108 44166
rect 27172 44102 27173 44166
rect 27659 44104 27660 44168
rect 27724 44104 27725 44168
rect 27659 44103 27725 44104
rect 27107 44101 27173 44102
rect 2099 43728 2165 43729
rect 2099 43726 2100 43728
rect 800 43666 2100 43726
rect 800 18042 1200 43666
rect 2099 43664 2100 43666
rect 2164 43664 2165 43728
rect 2099 43663 2165 43664
rect 800 18041 3498 18042
rect 800 17643 3099 18041
rect 3497 17643 3498 18041
rect 800 17642 3498 17643
rect 800 1000 1200 17642
rect 26498 1059 26678 1060
rect 26498 881 26499 1059
rect 26677 881 26678 1059
rect 3314 0 3494 200
rect 7178 0 7358 200
rect 11042 0 11222 200
rect 14906 0 15086 200
rect 18770 0 18950 200
rect 22634 0 22814 200
rect 26498 0 26678 881
rect 30362 921 30542 922
rect 30362 743 30363 921
rect 30541 743 30542 921
rect 30362 0 30542 743
use alt  alt_0
timestamp 1762479088
transform 1 0 18204 0 1 19994
box -3708 -3142 4491 1400
<< labels >>
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 29318 44952 29378 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 28214 44952 28274 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 30362 0 30542 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26498 0 26678 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22634 0 22814 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18770 0 18950 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 14906 0 15086 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 11042 0 11222 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 7178 0 7358 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 3314 0 3494 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 27662 44952 27722 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 27110 44952 27170 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 26006 44952 26066 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 25454 44952 25514 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 24902 44952 24962 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 23798 44952 23858 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23246 44952 23306 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22694 44952 22754 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21038 44952 21098 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 20486 44952 20546 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 19382 44952 19442 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 9998 44952 10058 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 9446 44952 9506 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 8342 44952 8402 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 7790 44952 7850 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 7238 44952 7298 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 6134 44952 6194 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 14414 44952 14474 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 13862 44952 13922 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 12758 44952 12818 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 12206 44952 12266 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 11654 44952 11714 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 10550 44952 10610 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 18830 44952 18890 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 18278 44952 18338 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 17174 44952 17234 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 16622 44952 16682 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 16070 44952 16130 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 14966 44952 15026 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 600 44152 1 FreeSans 400 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 800 1000 1200 44152 1 FreeSans 400 0 0 0 VGND
port 52 nsew ground bidirectional
flabel metal4 s 21590 44952 21650 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
