VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_analog_example
  CLASS BLOCK ;
  FOREIGN tt_um_analog_example ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 146.590 224.760 146.890 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 141.070 224.760 141.370 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 5.940000 ;
    ANTENNADIFFAREA 5.724000 ;
    PORT
      LAYER met4 ;
        RECT 151.810 0.000 152.710 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 5.940000 ;
    ANTENNADIFFAREA 5.724000 ;
    PORT
      LAYER met4 ;
        RECT 132.490 0.000 133.390 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 113.170 0.000 114.070 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 93.850 0.000 94.750 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 74.530 0.000 75.430 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.210 0.000 56.110 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 35.890 0.000 36.790 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 16.570 0.000 17.470 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 138.310 224.760 138.610 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 135.550 224.760 135.850 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 130.030 224.760 130.330 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 127.270 224.760 127.570 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 124.510 224.760 124.810 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.990 224.760 119.290 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 116.230 224.760 116.530 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 113.470 224.760 113.770 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.980000 ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.980000 ;
    PORT
      LAYER met4 ;
        RECT 107.950 224.760 108.250 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 105.190 224.760 105.490 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 102.430 224.760 102.730 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 96.910 224.760 97.210 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 49.990 224.760 50.290 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 47.230 224.760 47.530 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 41.710 224.760 42.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 38.950 224.760 39.250 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 36.190 224.760 36.490 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 30.670 224.760 30.970 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 72.070 224.760 72.370 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 69.310 224.760 69.610 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 63.790 224.760 64.090 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 61.030 224.760 61.330 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 58.270 224.760 58.570 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 52.750 224.760 53.050 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 94.150 224.760 94.450 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 91.390 224.760 91.690 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 85.870 224.760 86.170 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 83.110 224.760 83.410 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 80.350 224.760 80.650 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 74.830 224.760 75.130 225.760 ;
    END
  END uo_out[7]
  PIN VDPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 3.000 220.760 ;
    END
  END VDPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 4.000 5.000 6.000 220.760 ;
    END
  END VGND
  OBS
      LAYER pwell ;
        RECT 92.130 128.265 92.915 128.695 ;
        RECT 92.395 126.395 92.825 128.265 ;
      LAYER nwell ;
        RECT 93.245 128.060 94.850 128.900 ;
      LAYER pwell ;
        RECT 88.455 125.965 92.825 126.395 ;
        RECT 88.465 123.185 88.875 125.965 ;
      LAYER nwell ;
        RECT 93.710 125.560 94.550 128.060 ;
        RECT 89.180 123.955 96.920 125.560 ;
      LAYER pwell ;
        RECT 89.375 123.185 96.725 123.665 ;
        RECT 88.465 122.775 96.725 123.185 ;
        RECT 89.375 122.755 96.725 122.775 ;
        RECT 89.520 122.565 89.690 122.755 ;
        RECT 100.450 122.005 101.235 122.435 ;
        RECT 100.810 120.790 101.230 122.005 ;
      LAYER nwell ;
        RECT 101.565 121.800 103.170 122.640 ;
      LAYER pwell ;
        RECT 97.440 120.370 101.230 120.790 ;
      LAYER nwell ;
        RECT 87.690 118.065 97.080 119.670 ;
      LAYER pwell ;
        RECT 87.885 116.865 95.235 117.775 ;
        RECT 87.885 116.805 88.795 116.865 ;
        RECT 87.885 115.895 90.975 116.805 ;
      LAYER nwell ;
        RECT 95.475 116.125 97.080 118.065 ;
      LAYER pwell ;
        RECT 97.440 117.470 97.860 120.370 ;
      LAYER nwell ;
        RECT 101.920 119.730 102.760 121.800 ;
      LAYER pwell ;
        RECT 104.745 121.635 109.665 122.545 ;
      LAYER nwell ;
        RECT 109.995 121.800 111.600 122.640 ;
        RECT 98.510 118.125 103.030 119.730 ;
      LAYER pwell ;
        RECT 98.870 117.470 102.740 117.835 ;
        RECT 97.440 117.050 102.740 117.470 ;
        RECT 98.870 116.925 102.740 117.050 ;
        RECT 104.745 117.555 105.655 121.635 ;
      LAYER nwell ;
        RECT 110.380 119.450 111.220 121.800 ;
        RECT 106.290 117.845 114.030 119.450 ;
        RECT 116.500 117.775 124.620 119.380 ;
      LAYER pwell ;
        RECT 98.870 116.905 99.015 116.925 ;
        RECT 98.845 116.735 99.015 116.905 ;
        RECT 104.745 116.645 113.735 117.555 ;
        RECT 116.695 117.275 121.825 117.485 ;
        RECT 123.985 117.275 124.415 117.445 ;
        RECT 116.695 116.845 124.415 117.275 ;
        RECT 106.625 116.455 106.795 116.645 ;
        RECT 116.695 116.575 121.825 116.845 ;
        RECT 123.985 116.660 124.415 116.845 ;
        RECT 116.840 116.385 117.010 116.575 ;
        RECT 90.065 115.365 90.975 115.895 ;
      LAYER nwell ;
        RECT 92.380 115.570 97.080 116.125 ;
      LAYER pwell ;
        RECT 90.065 114.945 91.045 115.365 ;
        RECT 90.260 114.935 91.045 114.945 ;
      LAYER nwell ;
        RECT 91.375 114.730 97.080 115.570 ;
        RECT 92.380 114.520 97.080 114.730 ;
        RECT 95.475 114.470 97.080 114.520 ;
      LAYER pwell ;
        RECT 107.430 113.445 108.215 113.875 ;
        RECT 107.695 113.250 108.110 113.445 ;
        RECT 104.945 112.835 108.110 113.250 ;
      LAYER nwell ;
        RECT 108.545 113.240 110.150 114.080 ;
        RECT 82.180 111.570 83.020 111.740 ;
        RECT 82.180 110.135 95.710 111.570 ;
        RECT 82.800 109.965 95.710 110.135 ;
        RECT 98.400 109.955 104.470 111.560 ;
      LAYER pwell ;
        RECT 82.385 109.675 82.815 109.805 ;
        RECT 82.385 109.020 95.515 109.675 ;
        RECT 98.760 109.245 102.630 109.665 ;
        RECT 82.445 108.765 95.515 109.020 ;
        RECT 97.865 108.815 102.630 109.245 ;
        RECT 88.310 108.575 88.480 108.765 ;
        RECT 97.865 108.185 98.295 108.815 ;
        RECT 98.760 108.755 102.630 108.815 ;
        RECT 98.760 108.735 98.905 108.755 ;
        RECT 98.735 108.565 98.905 108.735 ;
        RECT 97.865 107.755 101.245 108.185 ;
        RECT 100.815 107.515 101.245 107.755 ;
      LAYER nwell ;
        RECT 102.865 107.720 104.470 109.955 ;
      LAYER pwell ;
        RECT 104.945 109.360 105.360 112.835 ;
      LAYER nwell ;
        RECT 108.910 111.560 109.750 113.240 ;
        RECT 106.290 109.955 114.030 111.560 ;
        RECT 116.250 111.390 124.470 111.430 ;
        RECT 116.250 109.825 125.100 111.390 ;
        RECT 124.260 109.785 125.100 109.825 ;
      LAYER pwell ;
        RECT 106.485 109.360 113.735 109.665 ;
        RECT 104.945 108.945 113.735 109.360 ;
        RECT 106.485 108.755 113.735 108.945 ;
        RECT 106.625 108.565 106.795 108.755 ;
        RECT 116.445 108.625 124.895 109.535 ;
        RECT 116.590 108.435 116.760 108.625 ;
        RECT 100.460 107.085 101.245 107.515 ;
      LAYER nwell ;
        RECT 101.575 106.880 104.470 107.720 ;
        RECT 102.865 106.850 104.470 106.880 ;
        RECT 99.440 105.910 100.280 106.140 ;
        RECT 88.860 104.535 100.280 105.910 ;
        RECT 88.860 104.305 99.840 104.535 ;
      LAYER pwell ;
        RECT 99.645 104.015 100.075 104.205 ;
        RECT 89.055 103.420 100.075 104.015 ;
        RECT 89.055 103.105 100.045 103.420 ;
        RECT 89.200 102.915 89.370 103.105 ;
      LAYER li1 ;
        RECT 91.855 128.625 92.025 128.710 ;
        RECT 94.575 128.625 94.745 128.710 ;
        RECT 91.855 128.335 92.750 128.625 ;
        RECT 93.410 128.335 94.745 128.625 ;
        RECT 91.855 128.250 92.025 128.335 ;
        RECT 94.575 128.250 94.745 128.335 ;
        RECT 89.370 125.285 96.730 125.455 ;
        RECT 89.460 124.145 89.715 125.285 ;
        RECT 89.885 124.315 90.215 125.115 ;
        RECT 90.385 124.485 90.555 125.285 ;
        RECT 90.725 124.315 91.055 125.115 ;
        RECT 91.225 124.485 91.395 125.285 ;
        RECT 91.565 124.315 91.895 125.115 ;
        RECT 92.065 124.485 92.235 125.285 ;
        RECT 92.405 124.315 92.735 125.115 ;
        RECT 92.905 124.485 93.075 125.285 ;
        RECT 93.245 124.315 93.575 125.115 ;
        RECT 93.745 124.485 93.915 125.285 ;
        RECT 94.085 124.315 94.415 125.115 ;
        RECT 94.585 124.485 94.755 125.285 ;
        RECT 94.925 124.315 95.255 125.115 ;
        RECT 95.425 124.485 95.595 125.285 ;
        RECT 95.765 124.315 96.095 125.115 ;
        RECT 89.885 124.115 96.095 124.315 ;
        RECT 96.285 124.145 96.640 125.285 ;
        RECT 89.880 123.725 92.735 123.945 ;
        RECT 93.010 123.725 93.490 124.115 ;
        RECT 93.660 123.725 95.675 123.925 ;
        RECT 93.245 123.555 93.490 123.725 ;
        RECT 95.845 123.555 96.095 124.115 ;
        RECT 89.460 123.385 93.075 123.555 ;
        RECT 89.460 122.905 89.795 123.385 ;
        RECT 89.965 122.735 90.135 123.215 ;
        RECT 90.305 122.905 90.635 123.385 ;
        RECT 90.805 122.735 90.975 123.215 ;
        RECT 91.145 122.905 91.475 123.385 ;
        RECT 91.645 122.735 91.815 123.215 ;
        RECT 91.985 122.905 92.315 123.385 ;
        RECT 92.485 122.735 92.655 123.215 ;
        RECT 92.825 123.135 93.075 123.385 ;
        RECT 93.245 123.305 96.095 123.555 ;
        RECT 96.265 123.135 96.640 123.555 ;
        RECT 92.825 122.905 96.640 123.135 ;
        RECT 89.370 122.565 96.730 122.735 ;
        RECT 100.175 122.365 100.345 122.450 ;
        RECT 102.895 122.365 103.065 122.450 ;
        RECT 100.175 122.075 101.070 122.365 ;
        RECT 101.730 122.075 103.065 122.365 ;
        RECT 100.175 121.990 100.345 122.075 ;
        RECT 102.895 121.990 103.065 122.075 ;
        RECT 108.605 122.365 108.775 122.450 ;
        RECT 111.325 122.365 111.495 122.450 ;
        RECT 108.605 122.075 109.500 122.365 ;
        RECT 110.160 122.075 111.495 122.365 ;
        RECT 108.605 121.990 108.775 122.075 ;
        RECT 111.325 121.990 111.495 122.075 ;
        RECT 87.880 119.395 95.240 119.565 ;
        RECT 98.700 119.455 102.840 119.625 ;
        RECT 87.970 118.255 88.225 119.395 ;
        RECT 88.395 118.425 88.725 119.225 ;
        RECT 88.895 118.595 89.065 119.395 ;
        RECT 89.235 118.425 89.565 119.225 ;
        RECT 89.735 118.595 89.905 119.395 ;
        RECT 90.075 118.425 90.405 119.225 ;
        RECT 90.575 118.595 90.745 119.395 ;
        RECT 90.915 118.425 91.245 119.225 ;
        RECT 91.415 118.595 91.585 119.395 ;
        RECT 91.755 118.425 92.085 119.225 ;
        RECT 92.255 118.595 92.425 119.395 ;
        RECT 92.595 118.425 92.925 119.225 ;
        RECT 93.095 118.595 93.265 119.395 ;
        RECT 93.435 118.425 93.765 119.225 ;
        RECT 93.935 118.595 94.105 119.395 ;
        RECT 94.275 118.425 94.605 119.225 ;
        RECT 88.395 118.225 94.605 118.425 ;
        RECT 94.795 118.255 95.150 119.395 ;
        RECT 98.955 118.655 99.210 119.455 ;
        RECT 99.380 118.485 99.710 119.285 ;
        RECT 99.880 118.655 100.050 119.455 ;
        RECT 100.220 118.485 100.550 119.285 ;
        RECT 100.720 118.655 100.890 119.455 ;
        RECT 101.060 118.485 101.390 119.285 ;
        RECT 101.560 118.655 101.730 119.455 ;
        RECT 101.900 118.485 102.230 119.285 ;
        RECT 102.400 118.655 102.700 119.455 ;
        RECT 106.480 119.175 113.840 119.345 ;
        RECT 98.785 118.315 102.755 118.485 ;
        RECT 88.390 117.835 91.245 118.055 ;
        RECT 91.520 117.835 92.000 118.225 ;
        RECT 92.170 117.835 94.185 118.035 ;
        RECT 91.755 117.665 92.000 117.835 ;
        RECT 94.355 117.665 94.605 118.225 ;
        RECT 98.785 117.725 99.130 118.315 ;
        RECT 99.380 117.895 102.235 118.145 ;
        RECT 102.435 117.725 102.755 118.315 ;
        RECT 106.570 118.205 106.885 119.005 ;
        RECT 107.055 118.375 107.305 119.175 ;
        RECT 107.475 118.205 107.725 119.005 ;
        RECT 107.895 118.375 108.145 119.175 ;
        RECT 108.315 118.205 108.565 119.005 ;
        RECT 108.735 118.375 108.985 119.175 ;
        RECT 109.155 118.205 109.405 119.005 ;
        RECT 109.575 118.375 109.825 119.175 ;
        RECT 116.690 119.105 122.210 119.275 ;
        RECT 123.970 119.105 124.430 119.275 ;
        RECT 109.995 118.835 113.605 119.005 ;
        RECT 109.995 118.205 110.245 118.835 ;
        RECT 106.570 117.995 110.245 118.205 ;
        RECT 110.415 118.155 110.665 118.665 ;
        RECT 110.835 118.325 111.085 118.835 ;
        RECT 111.255 118.155 111.505 118.665 ;
        RECT 111.675 118.325 111.925 118.835 ;
        RECT 112.095 118.155 112.345 118.665 ;
        RECT 112.515 118.325 112.765 118.835 ;
        RECT 112.935 118.155 113.185 118.665 ;
        RECT 113.355 118.325 113.605 118.835 ;
        RECT 110.415 117.985 113.755 118.155 ;
        RECT 87.970 117.495 91.585 117.665 ;
        RECT 87.970 117.015 88.305 117.495 ;
        RECT 88.475 116.845 88.645 117.325 ;
        RECT 88.815 117.015 89.145 117.495 ;
        RECT 89.315 116.845 89.485 117.325 ;
        RECT 89.655 117.015 89.985 117.495 ;
        RECT 90.155 116.845 90.325 117.325 ;
        RECT 90.495 117.015 90.825 117.495 ;
        RECT 90.995 116.845 91.165 117.325 ;
        RECT 91.335 117.245 91.585 117.495 ;
        RECT 91.755 117.415 94.605 117.665 ;
        RECT 94.775 117.245 95.150 117.665 ;
        RECT 98.785 117.535 102.755 117.725 ;
        RECT 106.840 117.615 110.010 117.815 ;
        RECT 110.280 117.615 113.020 117.815 ;
        RECT 91.335 117.015 95.150 117.245 ;
        RECT 98.955 116.905 99.210 117.365 ;
        RECT 99.380 117.075 99.710 117.535 ;
        RECT 99.880 116.905 100.050 117.365 ;
        RECT 100.220 117.075 100.550 117.535 ;
        RECT 100.720 116.905 100.890 117.365 ;
        RECT 101.060 117.075 101.390 117.535 ;
        RECT 101.560 116.905 101.730 117.365 ;
        RECT 101.900 117.075 102.230 117.535 ;
        RECT 113.190 117.445 113.755 117.985 ;
        RECT 116.785 118.085 117.115 118.935 ;
        RECT 117.285 118.305 117.455 119.105 ;
        RECT 117.625 118.085 117.955 118.935 ;
        RECT 118.125 118.305 118.295 119.105 ;
        RECT 118.545 118.085 118.715 118.935 ;
        RECT 118.885 118.305 119.215 119.105 ;
        RECT 119.385 118.085 119.555 118.935 ;
        RECT 119.725 118.305 120.055 119.105 ;
        RECT 120.225 118.085 120.395 118.935 ;
        RECT 120.565 118.305 120.895 119.105 ;
        RECT 121.065 118.085 121.235 118.935 ;
        RECT 116.785 117.915 118.285 118.085 ;
        RECT 118.545 117.915 121.235 118.085 ;
        RECT 121.405 117.955 121.735 119.105 ;
        RECT 124.055 117.940 124.345 119.105 ;
        RECT 116.830 117.545 117.930 117.745 ;
        RECT 118.110 117.715 118.285 117.915 ;
        RECT 118.110 117.545 120.735 117.715 ;
        RECT 102.400 116.905 102.705 117.365 ;
        RECT 87.880 116.675 95.240 116.845 ;
        RECT 98.700 116.735 102.840 116.905 ;
        RECT 106.570 116.625 106.845 117.445 ;
        RECT 107.015 117.265 113.755 117.445 ;
        RECT 118.110 117.375 118.285 117.545 ;
        RECT 120.980 117.375 121.235 117.915 ;
        RECT 107.015 116.795 107.345 117.265 ;
        RECT 107.515 116.625 107.685 117.095 ;
        RECT 107.855 116.795 108.185 117.265 ;
        RECT 108.355 116.625 108.525 117.095 ;
        RECT 108.695 116.795 109.025 117.265 ;
        RECT 109.195 116.625 109.365 117.095 ;
        RECT 109.535 116.795 109.865 117.265 ;
        RECT 110.035 116.625 110.205 117.095 ;
        RECT 110.375 116.795 110.705 117.265 ;
        RECT 110.875 116.625 111.045 117.095 ;
        RECT 111.215 116.795 111.545 117.265 ;
        RECT 111.715 116.625 111.885 117.095 ;
        RECT 112.055 116.795 112.385 117.265 ;
        RECT 112.555 116.625 112.725 117.095 ;
        RECT 112.895 116.795 113.225 117.265 ;
        RECT 116.865 117.205 118.285 117.375 ;
        RECT 118.545 117.205 121.235 117.375 ;
        RECT 113.395 116.625 113.685 117.095 ;
        RECT 116.865 116.725 117.035 117.205 ;
        RECT 106.480 116.455 113.840 116.625 ;
        RECT 117.205 116.555 117.535 117.035 ;
        RECT 117.705 116.730 117.875 117.205 ;
        RECT 118.045 116.555 118.375 117.035 ;
        RECT 118.545 116.725 118.715 117.205 ;
        RECT 118.885 116.555 119.215 117.035 ;
        RECT 119.385 116.725 119.555 117.205 ;
        RECT 119.725 116.555 120.055 117.035 ;
        RECT 120.225 116.725 120.395 117.205 ;
        RECT 120.565 116.555 120.895 117.035 ;
        RECT 121.065 116.725 121.235 117.205 ;
        RECT 121.405 116.555 121.735 117.355 ;
        RECT 124.055 116.555 124.345 117.280 ;
        RECT 116.690 116.385 122.210 116.555 ;
        RECT 123.970 116.385 124.430 116.555 ;
        RECT 89.985 115.295 90.155 115.380 ;
        RECT 92.705 115.295 92.875 115.380 ;
        RECT 89.985 115.005 90.880 115.295 ;
        RECT 91.540 115.005 92.875 115.295 ;
        RECT 89.985 114.920 90.155 115.005 ;
        RECT 92.705 114.920 92.875 115.005 ;
        RECT 107.155 113.805 107.325 113.890 ;
        RECT 109.875 113.805 110.045 113.890 ;
        RECT 107.155 113.515 108.050 113.805 ;
        RECT 108.710 113.515 110.045 113.805 ;
        RECT 107.155 113.430 107.325 113.515 ;
        RECT 109.875 113.430 110.045 113.515 ;
        RECT 82.370 111.465 82.830 111.635 ;
        RECT 82.455 110.300 82.745 111.465 ;
        RECT 88.160 111.295 95.520 111.465 ;
        RECT 88.250 110.155 88.505 111.295 ;
        RECT 88.675 110.325 89.005 111.125 ;
        RECT 89.175 110.495 89.345 111.295 ;
        RECT 89.515 110.325 89.845 111.125 ;
        RECT 90.015 110.495 90.185 111.295 ;
        RECT 90.355 110.325 90.685 111.125 ;
        RECT 90.855 110.495 91.025 111.295 ;
        RECT 91.195 110.325 91.525 111.125 ;
        RECT 91.695 110.495 91.865 111.295 ;
        RECT 92.035 110.325 92.365 111.125 ;
        RECT 92.535 110.495 92.705 111.295 ;
        RECT 92.875 110.325 93.205 111.125 ;
        RECT 93.375 110.495 93.545 111.295 ;
        RECT 93.715 110.325 94.045 111.125 ;
        RECT 94.215 110.495 94.385 111.295 ;
        RECT 94.555 110.325 94.885 111.125 ;
        RECT 88.675 110.125 94.885 110.325 ;
        RECT 95.075 110.155 95.430 111.295 ;
        RECT 98.590 111.285 102.730 111.455 ;
        RECT 106.480 111.285 113.840 111.455 ;
        RECT 98.845 110.485 99.100 111.285 ;
        RECT 99.270 110.315 99.600 111.115 ;
        RECT 99.770 110.485 99.940 111.285 ;
        RECT 100.110 110.315 100.440 111.115 ;
        RECT 100.610 110.485 100.780 111.285 ;
        RECT 100.950 110.315 101.280 111.115 ;
        RECT 101.450 110.485 101.620 111.285 ;
        RECT 101.790 110.315 102.120 111.115 ;
        RECT 102.290 110.485 102.590 111.285 ;
        RECT 106.570 110.315 106.885 111.115 ;
        RECT 107.055 110.485 107.305 111.285 ;
        RECT 107.475 110.315 107.725 111.115 ;
        RECT 107.895 110.485 108.145 111.285 ;
        RECT 108.315 110.315 108.565 111.115 ;
        RECT 108.735 110.485 108.985 111.285 ;
        RECT 109.155 110.315 109.405 111.115 ;
        RECT 109.575 110.485 109.825 111.285 ;
        RECT 116.440 111.155 121.960 111.325 ;
        RECT 109.995 110.945 113.605 111.115 ;
        RECT 109.995 110.315 110.245 110.945 ;
        RECT 88.670 109.735 91.525 109.955 ;
        RECT 91.800 109.735 92.280 110.125 ;
        RECT 92.450 109.735 94.465 109.935 ;
        RECT 82.455 108.915 82.745 109.640 ;
        RECT 92.035 109.565 92.280 109.735 ;
        RECT 94.635 109.565 94.885 110.125 ;
        RECT 98.675 110.145 102.645 110.315 ;
        RECT 88.250 109.395 91.865 109.565 ;
        RECT 88.250 108.915 88.585 109.395 ;
        RECT 82.370 108.745 82.830 108.915 ;
        RECT 88.755 108.745 88.925 109.225 ;
        RECT 89.095 108.915 89.425 109.395 ;
        RECT 89.595 108.745 89.765 109.225 ;
        RECT 89.935 108.915 90.265 109.395 ;
        RECT 90.435 108.745 90.605 109.225 ;
        RECT 90.775 108.915 91.105 109.395 ;
        RECT 91.275 108.745 91.445 109.225 ;
        RECT 91.615 109.145 91.865 109.395 ;
        RECT 92.035 109.315 94.885 109.565 ;
        RECT 95.055 109.145 95.430 109.565 ;
        RECT 98.675 109.555 99.020 110.145 ;
        RECT 99.270 109.725 102.125 109.975 ;
        RECT 102.325 109.555 102.645 110.145 ;
        RECT 106.570 110.105 110.245 110.315 ;
        RECT 110.415 110.265 110.665 110.775 ;
        RECT 110.835 110.435 111.085 110.945 ;
        RECT 111.255 110.265 111.505 110.775 ;
        RECT 111.675 110.435 111.925 110.945 ;
        RECT 112.095 110.265 112.345 110.775 ;
        RECT 112.515 110.435 112.765 110.945 ;
        RECT 112.935 110.265 113.185 110.775 ;
        RECT 113.355 110.435 113.605 110.945 ;
        RECT 110.415 110.095 113.755 110.265 ;
        RECT 106.840 109.725 110.010 109.925 ;
        RECT 110.280 109.725 113.020 109.925 ;
        RECT 113.190 109.555 113.755 110.095 ;
        RECT 116.535 110.135 116.865 110.985 ;
        RECT 117.035 110.355 117.205 111.155 ;
        RECT 117.375 110.135 117.705 110.985 ;
        RECT 117.875 110.355 118.045 111.155 ;
        RECT 118.295 110.135 118.465 110.985 ;
        RECT 118.635 110.355 118.965 111.155 ;
        RECT 119.135 110.135 119.305 110.985 ;
        RECT 119.475 110.355 119.805 111.155 ;
        RECT 119.975 110.135 120.145 110.985 ;
        RECT 120.315 110.355 120.645 111.155 ;
        RECT 120.815 110.135 120.985 110.985 ;
        RECT 116.535 109.965 118.035 110.135 ;
        RECT 118.295 109.965 120.985 110.135 ;
        RECT 121.155 110.005 121.485 111.155 ;
        RECT 124.450 111.115 124.910 111.285 ;
        RECT 116.580 109.595 117.680 109.795 ;
        RECT 117.860 109.765 118.035 109.965 ;
        RECT 117.860 109.595 120.485 109.765 ;
        RECT 98.675 109.365 102.645 109.555 ;
        RECT 91.615 108.915 95.430 109.145 ;
        RECT 88.160 108.575 95.520 108.745 ;
        RECT 98.845 108.735 99.100 109.195 ;
        RECT 99.270 108.905 99.600 109.365 ;
        RECT 99.770 108.735 99.940 109.195 ;
        RECT 100.110 108.905 100.440 109.365 ;
        RECT 100.610 108.735 100.780 109.195 ;
        RECT 100.950 108.905 101.280 109.365 ;
        RECT 101.450 108.735 101.620 109.195 ;
        RECT 101.790 108.905 102.120 109.365 ;
        RECT 102.290 108.735 102.595 109.195 ;
        RECT 106.570 108.735 106.845 109.555 ;
        RECT 107.015 109.375 113.755 109.555 ;
        RECT 117.860 109.425 118.035 109.595 ;
        RECT 120.730 109.425 120.985 109.965 ;
        RECT 124.535 109.950 124.825 111.115 ;
        RECT 107.015 108.905 107.345 109.375 ;
        RECT 107.515 108.735 107.685 109.205 ;
        RECT 107.855 108.905 108.185 109.375 ;
        RECT 108.355 108.735 108.525 109.205 ;
        RECT 108.695 108.905 109.025 109.375 ;
        RECT 109.195 108.735 109.365 109.205 ;
        RECT 109.535 108.905 109.865 109.375 ;
        RECT 110.035 108.735 110.205 109.205 ;
        RECT 110.375 108.905 110.705 109.375 ;
        RECT 110.875 108.735 111.045 109.205 ;
        RECT 111.215 108.905 111.545 109.375 ;
        RECT 111.715 108.735 111.885 109.205 ;
        RECT 112.055 108.905 112.385 109.375 ;
        RECT 112.555 108.735 112.725 109.205 ;
        RECT 112.895 108.905 113.225 109.375 ;
        RECT 116.615 109.255 118.035 109.425 ;
        RECT 118.295 109.255 120.985 109.425 ;
        RECT 113.395 108.735 113.685 109.205 ;
        RECT 116.615 108.775 116.785 109.255 ;
        RECT 98.590 108.565 102.730 108.735 ;
        RECT 106.480 108.565 113.840 108.735 ;
        RECT 116.955 108.605 117.285 109.085 ;
        RECT 117.455 108.780 117.625 109.255 ;
        RECT 117.795 108.605 118.125 109.085 ;
        RECT 118.295 108.775 118.465 109.255 ;
        RECT 118.635 108.605 118.965 109.085 ;
        RECT 119.135 108.775 119.305 109.255 ;
        RECT 119.475 108.605 119.805 109.085 ;
        RECT 119.975 108.775 120.145 109.255 ;
        RECT 120.315 108.605 120.645 109.085 ;
        RECT 120.815 108.775 120.985 109.255 ;
        RECT 121.155 108.605 121.485 109.405 ;
        RECT 116.440 108.435 121.960 108.605 ;
        RECT 124.535 108.565 124.825 109.290 ;
        RECT 124.450 108.395 124.910 108.565 ;
        RECT 100.185 107.445 100.355 107.530 ;
        RECT 102.905 107.445 103.075 107.530 ;
        RECT 100.185 107.155 101.080 107.445 ;
        RECT 101.740 107.155 103.075 107.445 ;
        RECT 100.185 107.070 100.355 107.155 ;
        RECT 102.905 107.070 103.075 107.155 ;
        RECT 99.630 105.865 100.090 106.035 ;
        RECT 89.050 105.635 96.410 105.805 ;
        RECT 89.140 104.495 89.395 105.635 ;
        RECT 89.565 104.665 89.895 105.465 ;
        RECT 90.065 104.835 90.235 105.635 ;
        RECT 90.405 104.665 90.735 105.465 ;
        RECT 90.905 104.835 91.075 105.635 ;
        RECT 91.245 104.665 91.575 105.465 ;
        RECT 91.745 104.835 91.915 105.635 ;
        RECT 92.085 104.665 92.415 105.465 ;
        RECT 92.585 104.835 92.755 105.635 ;
        RECT 92.925 104.665 93.255 105.465 ;
        RECT 93.425 104.835 93.595 105.635 ;
        RECT 93.765 104.665 94.095 105.465 ;
        RECT 94.265 104.835 94.435 105.635 ;
        RECT 94.605 104.665 94.935 105.465 ;
        RECT 95.105 104.835 95.275 105.635 ;
        RECT 95.445 104.665 95.775 105.465 ;
        RECT 89.565 104.465 95.775 104.665 ;
        RECT 95.965 104.495 96.320 105.635 ;
        RECT 99.715 104.700 100.005 105.865 ;
        RECT 89.560 104.075 92.415 104.295 ;
        RECT 92.690 104.075 93.170 104.465 ;
        RECT 93.340 104.075 95.355 104.275 ;
        RECT 92.925 103.905 93.170 104.075 ;
        RECT 95.525 103.905 95.775 104.465 ;
        RECT 89.140 103.735 92.755 103.905 ;
        RECT 89.140 103.255 89.475 103.735 ;
        RECT 89.645 103.085 89.815 103.565 ;
        RECT 89.985 103.255 90.315 103.735 ;
        RECT 90.485 103.085 90.655 103.565 ;
        RECT 90.825 103.255 91.155 103.735 ;
        RECT 91.325 103.085 91.495 103.565 ;
        RECT 91.665 103.255 91.995 103.735 ;
        RECT 92.165 103.085 92.335 103.565 ;
        RECT 92.505 103.485 92.755 103.735 ;
        RECT 92.925 103.655 95.775 103.905 ;
        RECT 95.945 103.485 96.320 103.905 ;
        RECT 92.505 103.255 96.320 103.485 ;
        RECT 99.715 103.315 100.005 104.040 ;
        RECT 99.630 103.145 100.090 103.315 ;
        RECT 89.050 102.915 96.410 103.085 ;
      LAYER met1 ;
        RECT 113.440 147.560 113.800 147.860 ;
        RECT 113.470 136.615 113.770 147.560 ;
        RECT 128.470 139.620 128.730 139.940 ;
        RECT 112.635 136.360 127.015 136.615 ;
        RECT 85.900 136.030 86.160 136.350 ;
        RECT 85.920 123.945 86.140 136.030 ;
        RECT 91.700 128.250 92.180 128.710 ;
        RECT 94.420 128.250 94.900 128.710 ;
        RECT 91.700 126.735 91.855 128.250 ;
        RECT 91.620 126.475 91.940 126.735 ;
        RECT 87.135 125.610 87.425 125.640 ;
        RECT 94.745 125.610 94.900 128.250 ;
        RECT 87.135 125.455 103.985 125.610 ;
        RECT 87.135 125.320 96.730 125.455 ;
        RECT 87.135 125.290 87.425 125.320 ;
        RECT 89.370 125.130 96.730 125.320 ;
        RECT 92.840 124.210 93.690 124.310 ;
        RECT 90.130 123.945 90.410 123.975 ;
        RECT 85.920 123.725 90.800 123.945 ;
        RECT 92.840 123.830 99.030 124.210 ;
        RECT 100.680 124.070 100.980 124.100 ;
        RECT 92.850 123.730 99.030 123.830 ;
        RECT 92.890 123.725 99.030 123.730 ;
        RECT 90.130 123.695 90.410 123.725 ;
        RECT 92.890 123.470 93.690 123.725 ;
        RECT 95.160 123.665 95.420 123.725 ;
        RECT 89.370 122.625 96.730 122.890 ;
        RECT 86.275 122.470 96.730 122.625 ;
        RECT 86.275 119.720 86.430 122.470 ;
        RECT 89.370 122.410 96.730 122.470 ;
        RECT 90.195 121.935 90.350 122.410 ;
        RECT 90.140 121.615 90.400 121.935 ;
        RECT 98.550 121.220 99.030 123.725 ;
        RECT 100.040 123.770 100.980 124.070 ;
        RECT 100.040 122.450 100.340 123.770 ;
        RECT 100.680 123.740 100.980 123.770 ;
        RECT 100.020 121.990 100.500 122.450 ;
        RECT 102.740 121.990 103.220 122.450 ;
        RECT 96.860 120.740 99.030 121.220 ;
        RECT 93.460 119.720 93.760 120.090 ;
        RECT 86.270 119.565 86.440 119.720 ;
        RECT 87.880 119.635 95.240 119.720 ;
        RECT 86.275 116.675 86.430 119.565 ;
        RECT 87.105 119.345 95.240 119.635 ;
        RECT 87.880 119.240 95.240 119.345 ;
        RECT 95.900 118.820 96.440 119.300 ;
        RECT 91.490 118.315 92.030 118.345 ;
        RECT 89.040 118.055 89.320 118.085 ;
        RECT 87.100 117.835 89.770 118.055 ;
        RECT 91.230 117.835 92.160 118.315 ;
        RECT 96.005 118.295 96.340 118.820 ;
        RECT 96.860 118.295 97.340 120.740 ;
        RECT 98.700 119.630 102.840 119.780 ;
        RECT 103.065 119.630 103.220 121.990 ;
        RECT 103.830 119.630 103.985 125.455 ;
        RECT 104.935 122.180 105.195 122.265 ;
        RECT 108.450 122.180 108.930 122.450 ;
        RECT 104.935 122.025 108.930 122.180 ;
        RECT 104.935 121.945 105.195 122.025 ;
        RECT 108.450 121.990 108.930 122.025 ;
        RECT 111.170 121.990 111.650 122.450 ;
        RECT 98.700 119.500 105.595 119.630 ;
        RECT 111.495 119.500 111.650 121.990 ;
        RECT 98.700 119.475 113.840 119.500 ;
        RECT 98.700 119.300 102.840 119.475 ;
        RECT 105.440 119.430 113.840 119.475 ;
        RECT 105.440 119.345 124.430 119.430 ;
        RECT 105.440 119.340 105.595 119.345 ;
        RECT 106.480 119.275 124.430 119.345 ;
        RECT 106.480 119.020 113.840 119.275 ;
        RECT 116.690 118.950 122.210 119.275 ;
        RECT 123.970 118.950 124.430 119.275 ;
        RECT 96.000 118.145 97.340 118.295 ;
        RECT 100.020 118.145 100.330 118.175 ;
        RECT 93.690 118.035 93.950 118.065 ;
        RECT 95.010 118.035 95.330 118.065 ;
        RECT 93.390 117.835 95.330 118.035 ;
        RECT 87.100 117.510 87.320 117.835 ;
        RECT 89.040 117.805 89.320 117.835 ;
        RECT 91.490 117.805 92.030 117.835 ;
        RECT 93.690 117.805 93.950 117.835 ;
        RECT 95.010 117.805 95.330 117.835 ;
        RECT 96.000 117.895 100.505 118.145 ;
        RECT 102.405 118.120 102.785 118.150 ;
        RECT 102.160 117.930 105.830 118.120 ;
        RECT 113.160 117.955 113.785 118.015 ;
        RECT 114.640 117.960 115.205 118.660 ;
        RECT 114.590 117.955 115.205 117.960 ;
        RECT 96.000 117.890 97.340 117.895 ;
        RECT 96.000 117.855 97.330 117.890 ;
        RECT 100.020 117.865 100.330 117.895 ;
        RECT 96.000 117.730 96.290 117.855 ;
        RECT 102.160 117.800 107.490 117.930 ;
        RECT 102.405 117.770 102.785 117.800 ;
        RECT 105.500 117.785 107.490 117.800 ;
        RECT 109.175 117.785 109.405 117.815 ;
        RECT 87.080 117.190 87.340 117.510 ;
        RECT 95.990 117.310 96.290 117.730 ;
        RECT 105.500 117.615 109.675 117.785 ;
        RECT 105.500 117.610 107.490 117.615 ;
        RECT 109.175 117.585 109.405 117.615 ;
        RECT 110.615 117.525 111.225 117.895 ;
        RECT 113.160 117.745 115.880 117.955 ;
        RECT 117.075 117.745 117.325 117.805 ;
        RECT 113.160 117.555 117.325 117.745 ;
        RECT 110.615 117.515 111.005 117.525 ;
        RECT 113.160 117.390 115.880 117.555 ;
        RECT 117.075 117.495 117.325 117.555 ;
        RECT 120.950 117.710 121.265 117.770 ;
        RECT 126.760 117.710 127.015 136.360 ;
        RECT 120.950 117.455 127.015 117.710 ;
        RECT 120.950 117.390 121.265 117.455 ;
        RECT 113.160 117.320 113.785 117.390 ;
        RECT 95.960 117.010 96.320 117.310 ;
        RECT 87.880 116.675 95.240 117.000 ;
        RECT 98.110 116.825 98.370 116.910 ;
        RECT 98.700 116.825 102.840 117.060 ;
        RECT 97.505 116.735 102.840 116.825 ;
        RECT 97.505 116.675 105.475 116.735 ;
        RECT 86.275 116.525 97.655 116.675 ;
        RECT 98.110 116.590 98.370 116.675 ;
        RECT 98.700 116.580 105.475 116.675 ;
        RECT 86.275 116.520 95.240 116.525 ;
        RECT 82.755 115.485 83.105 115.775 ;
        RECT 41.515 115.275 55.550 115.450 ;
        RECT 41.515 115.165 69.935 115.275 ;
        RECT 82.785 115.165 83.075 115.485 ;
        RECT 88.265 115.270 88.420 116.520 ;
        RECT 105.320 116.500 105.475 116.580 ;
        RECT 106.480 116.500 113.840 116.780 ;
        RECT 114.590 116.770 115.155 117.390 ;
        RECT 105.320 116.455 113.840 116.500 ;
        RECT 115.355 116.455 115.510 116.460 ;
        RECT 116.690 116.455 122.210 116.710 ;
        RECT 105.320 116.385 122.210 116.455 ;
        RECT 123.970 116.385 124.430 116.710 ;
        RECT 105.320 116.345 124.430 116.385 ;
        RECT 106.480 116.300 124.430 116.345 ;
        RECT 89.830 115.270 90.310 115.380 ;
        RECT 41.515 114.875 83.075 115.165 ;
        RECT 41.515 114.765 69.935 114.875 ;
        RECT 41.515 114.595 55.550 114.765 ;
        RECT 82.785 112.295 83.075 114.875 ;
        RECT 85.475 115.115 90.310 115.270 ;
        RECT 85.475 113.435 85.630 115.115 ;
        RECT 89.830 114.920 90.310 115.115 ;
        RECT 92.550 115.305 93.030 115.380 ;
        RECT 93.650 115.305 93.970 115.360 ;
        RECT 107.140 115.350 107.440 116.300 ;
        RECT 115.355 116.270 115.510 116.300 ;
        RECT 116.690 116.230 124.430 116.300 ;
        RECT 92.550 115.150 93.970 115.305 ;
        RECT 114.560 115.240 115.185 115.805 ;
        RECT 92.550 114.920 93.030 115.150 ;
        RECT 93.650 115.100 93.970 115.150 ;
        RECT 114.590 115.015 115.155 115.240 ;
        RECT 103.130 114.450 115.155 115.015 ;
        RECT 107.000 113.690 107.480 113.890 ;
        RECT 105.035 113.535 107.480 113.690 ;
        RECT 85.425 113.115 85.685 113.435 ;
        RECT 105.035 112.995 105.190 113.535 ;
        RECT 107.000 113.430 107.480 113.535 ;
        RECT 109.720 113.430 110.200 113.890 ;
        RECT 104.985 112.675 105.245 112.995 ;
        RECT 110.045 112.925 110.200 113.430 ;
        RECT 82.655 112.140 88.805 112.295 ;
        RECT 82.655 112.125 83.075 112.140 ;
        RECT 82.655 111.790 82.810 112.125 ;
        RECT 82.370 111.310 82.830 111.790 ;
        RECT 88.650 111.620 88.805 112.140 ;
        RECT 88.160 111.610 98.825 111.620 ;
        RECT 100.860 111.610 101.160 112.640 ;
        RECT 109.995 112.605 110.255 112.925 ;
        RECT 110.450 112.215 110.770 112.260 ;
        RECT 105.535 112.045 110.770 112.215 ;
        RECT 105.535 111.790 105.705 112.045 ;
        RECT 110.450 112.000 110.770 112.045 ;
        RECT 105.535 111.705 105.715 111.790 ;
        RECT 104.370 111.610 104.690 111.665 ;
        RECT 88.160 111.465 104.690 111.610 ;
        RECT 87.130 111.400 87.450 111.450 ;
        RECT 88.160 111.400 95.520 111.465 ;
        RECT 87.130 111.245 95.520 111.400 ;
        RECT 87.130 111.190 87.450 111.245 ;
        RECT 88.160 111.140 95.520 111.245 ;
        RECT 98.590 111.455 104.690 111.465 ;
        RECT 98.590 111.130 102.730 111.455 ;
        RECT 104.370 111.405 104.690 111.455 ;
        RECT 91.800 110.245 92.280 110.520 ;
        RECT 96.060 110.330 96.320 110.650 ;
        RECT 90.185 109.955 90.465 110.015 ;
        RECT 84.560 109.735 90.465 109.955 ;
        RECT 82.370 108.745 82.830 109.070 ;
        RECT 83.190 108.745 83.510 108.800 ;
        RECT 82.370 108.590 83.510 108.745 ;
        RECT 83.190 108.540 83.510 108.590 ;
        RECT 84.560 102.620 84.780 109.735 ;
        RECT 90.185 109.675 90.465 109.735 ;
        RECT 91.770 109.705 92.310 110.245 ;
        RECT 93.980 109.935 94.240 109.965 ;
        RECT 96.090 109.935 96.290 110.330 ;
        RECT 93.800 109.735 96.290 109.935 ;
        RECT 99.170 109.975 99.490 109.980 ;
        RECT 99.910 109.975 100.220 110.005 ;
        RECT 102.295 109.980 102.675 110.010 ;
        RECT 93.980 109.705 94.240 109.735 ;
        RECT 99.170 109.725 100.785 109.975 ;
        RECT 102.180 109.885 104.240 109.980 ;
        RECT 105.545 109.885 105.715 111.705 ;
        RECT 109.970 111.610 110.290 111.855 ;
        RECT 105.980 111.385 106.240 111.465 ;
        RECT 106.480 111.455 115.355 111.610 ;
        RECT 106.480 111.385 113.840 111.455 ;
        RECT 105.980 111.230 113.840 111.385 ;
        RECT 105.980 111.145 106.240 111.230 ;
        RECT 106.480 111.130 113.840 111.230 ;
        RECT 115.200 111.370 115.355 111.455 ;
        RECT 116.440 111.440 121.960 111.480 ;
        RECT 116.440 111.370 124.910 111.440 ;
        RECT 115.200 111.285 124.910 111.370 ;
        RECT 115.200 111.215 121.960 111.285 ;
        RECT 116.440 111.000 121.960 111.215 ;
        RECT 124.450 110.960 124.910 111.285 ;
        RECT 115.280 110.420 115.540 110.740 ;
        RECT 113.160 110.270 113.785 110.325 ;
        RECT 110.540 110.005 110.710 110.035 ;
        RECT 107.475 109.895 107.705 109.925 ;
        RECT 99.170 109.720 99.490 109.725 ;
        RECT 91.800 109.390 92.280 109.705 ;
        RECT 99.910 109.695 100.220 109.725 ;
        RECT 102.180 109.715 105.715 109.885 ;
        RECT 106.075 109.725 107.935 109.895 ;
        RECT 102.180 109.660 104.240 109.715 ;
        RECT 102.295 109.630 102.675 109.660 ;
        RECT 105.370 109.285 105.690 109.330 ;
        RECT 106.075 109.285 106.245 109.725 ;
        RECT 107.475 109.695 107.705 109.725 ;
        RECT 110.445 109.655 110.885 110.005 ;
        RECT 113.160 109.775 114.800 110.270 ;
        RECT 115.325 109.775 115.495 110.420 ;
        RECT 120.715 109.850 120.970 109.945 ;
        RECT 120.700 109.820 121.015 109.850 ;
        RECT 116.800 109.775 117.030 109.805 ;
        RECT 120.595 109.785 121.965 109.820 ;
        RECT 128.485 109.785 128.715 139.620 ;
        RECT 113.160 109.705 117.305 109.775 ;
        RECT 110.445 109.635 110.785 109.655 ;
        RECT 113.160 109.640 113.785 109.705 ;
        RECT 110.480 109.560 110.740 109.635 ;
        RECT 114.235 109.605 117.305 109.705 ;
        RECT 87.155 108.800 87.415 109.120 ;
        RECT 105.370 109.115 106.245 109.285 ;
        RECT 105.370 109.070 105.690 109.115 ;
        RECT 87.205 105.960 87.360 108.800 ;
        RECT 88.160 108.660 95.520 108.900 ;
        RECT 97.835 108.660 97.990 108.665 ;
        RECT 98.590 108.660 102.730 108.890 ;
        RECT 106.480 108.660 113.840 108.890 ;
        RECT 88.160 108.565 113.840 108.660 ;
        RECT 88.160 108.505 114.025 108.565 ;
        RECT 88.160 108.420 95.520 108.505 ;
        RECT 88.970 107.600 89.270 108.420 ;
        RECT 96.770 107.300 97.250 108.040 ;
        RECT 97.835 107.325 97.990 108.505 ;
        RECT 98.590 108.410 102.730 108.505 ;
        RECT 106.480 108.410 114.025 108.505 ;
        RECT 103.025 107.820 103.285 108.140 ;
        RECT 103.075 107.530 103.230 107.820 ;
        RECT 100.030 107.325 100.510 107.530 ;
        RECT 96.785 106.900 97.195 107.300 ;
        RECT 97.835 107.170 100.510 107.325 ;
        RECT 96.750 106.360 97.230 106.900 ;
        RECT 96.860 106.070 97.060 106.360 ;
        RECT 87.205 105.805 96.410 105.960 ;
        RECT 96.860 105.870 97.510 106.070 ;
        RECT 89.050 105.695 96.410 105.805 ;
        RECT 89.050 105.540 96.885 105.695 ;
        RECT 89.050 105.480 96.410 105.540 ;
        RECT 96.730 105.180 96.885 105.540 ;
        RECT 96.645 104.920 96.965 105.180 ;
        RECT 92.660 104.555 93.200 104.585 ;
        RECT 85.700 104.295 86.020 104.315 ;
        RECT 90.205 104.295 90.485 104.325 ;
        RECT 85.700 104.075 91.000 104.295 ;
        RECT 92.410 104.075 93.350 104.555 ;
        RECT 94.875 104.275 95.135 104.305 ;
        RECT 97.310 104.275 97.510 105.870 ;
        RECT 94.240 104.075 97.510 104.275 ;
        RECT 85.700 104.055 86.020 104.075 ;
        RECT 90.205 104.045 90.485 104.075 ;
        RECT 92.660 104.045 93.200 104.075 ;
        RECT 94.875 104.045 95.135 104.075 ;
        RECT 89.050 103.110 96.410 103.240 ;
        RECT 97.835 103.185 97.990 107.170 ;
        RECT 100.030 107.070 100.510 107.170 ;
        RECT 102.750 107.070 103.230 107.530 ;
        RECT 106.640 107.780 106.940 107.810 ;
        RECT 107.240 107.780 107.540 108.410 ;
        RECT 113.870 108.005 114.025 108.410 ;
        RECT 106.640 107.480 107.540 107.780 ;
        RECT 113.820 107.685 114.080 108.005 ;
        RECT 106.640 107.450 106.940 107.480 ;
        RECT 114.235 107.060 114.800 109.605 ;
        RECT 116.800 109.575 117.030 109.605 ;
        RECT 120.595 109.565 128.715 109.785 ;
        RECT 120.700 109.555 128.715 109.565 ;
        RECT 120.700 109.530 121.285 109.555 ;
        RECT 120.715 109.365 121.285 109.530 ;
        RECT 116.440 108.520 121.960 108.760 ;
        RECT 124.450 108.520 124.910 108.720 ;
        RECT 116.440 108.420 124.910 108.520 ;
        RECT 115.870 108.375 124.910 108.420 ;
        RECT 115.870 108.280 121.960 108.375 ;
        RECT 115.870 108.200 116.630 108.280 ;
        RECT 124.450 108.240 124.910 108.375 ;
        RECT 115.870 108.005 116.090 108.200 ;
        RECT 115.850 107.685 116.110 108.005 ;
        RECT 110.390 106.840 114.850 107.060 ;
        RECT 98.935 106.035 100.090 106.190 ;
        RECT 98.935 105.205 99.090 106.035 ;
        RECT 99.630 105.710 100.090 106.035 ;
        RECT 98.885 104.885 99.145 105.205 ;
        RECT 99.630 103.185 100.090 103.470 ;
        RECT 97.835 103.110 100.090 103.185 ;
        RECT 89.050 102.990 100.090 103.110 ;
        RECT 89.050 102.955 99.845 102.990 ;
        RECT 89.050 102.760 96.410 102.955 ;
        RECT 110.390 102.620 110.610 106.840 ;
        RECT 112.450 106.780 114.800 106.840 ;
        RECT 84.560 102.400 110.610 102.620 ;
      LAYER met2 ;
        RECT 116.230 179.820 116.530 179.830 ;
        RECT 116.195 179.540 116.565 179.820 ;
        RECT 113.470 179.190 113.770 179.200 ;
        RECT 113.435 178.910 113.805 179.190 ;
        RECT 85.880 151.195 86.180 151.585 ;
        RECT 85.920 136.320 86.140 151.195 ;
        RECT 113.470 147.530 113.770 178.910 ;
        RECT 116.230 139.895 116.530 179.540 ;
        RECT 128.440 139.895 128.760 139.910 ;
        RECT 114.735 139.665 128.760 139.895 ;
        RECT 128.440 139.650 128.760 139.665 ;
        RECT 85.870 136.060 86.190 136.320 ;
        RECT 91.650 126.685 91.910 126.765 ;
        RECT 87.975 126.530 91.910 126.685 ;
        RECT 87.105 125.320 87.455 125.610 ;
        RECT 87.135 120.335 87.425 125.320 ;
        RECT 87.975 121.850 88.130 126.530 ;
        RECT 91.650 126.445 91.910 126.530 ;
        RECT 100.650 124.060 101.010 124.070 ;
        RECT 100.645 123.780 101.015 124.060 ;
        RECT 100.650 123.770 101.010 123.780 ;
        RECT 104.990 122.235 105.145 122.465 ;
        RECT 104.905 121.975 105.225 122.235 ;
        RECT 90.110 121.850 90.430 121.905 ;
        RECT 87.975 121.695 90.430 121.850 ;
        RECT 104.920 121.840 105.220 121.975 ;
        RECT 104.990 121.795 105.145 121.840 ;
        RECT 90.110 121.645 90.430 121.695 ;
        RECT 84.585 120.045 87.425 120.335 ;
        RECT 82.785 115.775 83.075 115.805 ;
        RECT 84.585 115.775 84.875 120.045 ;
        RECT 87.135 119.315 87.425 120.045 ;
        RECT 91.650 117.805 92.130 120.905 ;
        RECT 99.360 120.630 115.205 121.180 ;
        RECT 97.610 120.615 115.205 120.630 ;
        RECT 97.610 120.150 99.925 120.615 ;
        RECT 93.470 120.060 93.750 120.095 ;
        RECT 93.430 119.760 93.790 120.060 ;
        RECT 93.470 119.725 93.750 119.760 ;
        RECT 95.930 119.725 96.410 119.750 ;
        RECT 95.910 119.295 96.430 119.725 ;
        RECT 95.930 118.790 96.410 119.295 ;
        RECT 97.610 118.110 98.090 120.150 ;
        RECT 99.360 120.110 99.925 120.150 ;
        RECT 114.640 118.630 115.205 120.615 ;
        RECT 95.260 118.095 98.090 118.110 ;
        RECT 95.040 117.775 98.090 118.095 ;
        RECT 114.610 118.065 115.235 118.630 ;
        RECT 95.260 117.710 98.090 117.775 ;
        RECT 97.610 117.670 98.090 117.710 ;
        RECT 110.810 117.570 111.070 117.890 ;
        RECT 87.050 117.220 87.370 117.480 ;
        RECT 82.785 115.485 84.875 115.775 ;
        RECT 41.545 115.450 42.400 115.480 ;
        RECT 82.785 115.455 83.075 115.485 ;
        RECT 13.340 114.595 42.400 115.450 ;
        RECT 41.545 114.565 42.400 114.595 ;
        RECT 87.100 114.180 87.320 117.220 ;
        RECT 95.990 116.280 96.290 117.340 ;
        RECT 98.090 116.880 98.390 116.945 ;
        RECT 98.080 116.620 98.400 116.880 ;
        RECT 98.090 116.555 98.390 116.620 ;
        RECT 95.990 115.980 100.395 116.280 ;
        RECT 110.855 116.095 111.025 117.570 ;
        RECT 114.560 116.800 115.185 117.365 ;
        RECT 95.990 115.690 96.290 115.980 ;
        RECT 110.710 115.915 111.025 116.095 ;
        RECT 95.955 115.410 96.325 115.690 ;
        RECT 106.570 115.680 106.850 115.715 ;
        RECT 93.680 115.380 93.940 115.390 ;
        RECT 106.130 115.380 107.470 115.680 ;
        RECT 110.710 115.595 110.895 115.915 ;
        RECT 93.615 115.080 94.005 115.380 ;
        RECT 106.570 115.345 106.850 115.380 ;
        RECT 110.710 115.280 110.900 115.595 ;
        RECT 93.680 115.070 93.940 115.080 ;
        RECT 103.250 114.420 103.815 115.045 ;
        RECT 99.965 114.180 100.355 114.220 ;
        RECT 87.100 113.960 100.355 114.180 ;
        RECT 85.395 113.355 85.715 113.405 ;
        RECT 51.910 113.090 65.925 113.205 ;
        RECT 83.950 113.195 85.715 113.355 ;
        RECT 95.790 113.350 96.470 113.650 ;
        RECT 51.910 112.975 70.350 113.090 ;
        RECT 51.910 112.890 75.585 112.975 ;
        RECT 83.950 112.890 84.110 113.195 ;
        RECT 85.395 113.145 85.715 113.195 ;
        RECT 51.910 112.730 84.110 112.890 ;
        RECT 51.910 112.645 75.585 112.730 ;
        RECT 51.910 112.530 70.350 112.645 ;
        RECT 51.910 112.415 65.925 112.530 ;
        RECT 83.220 108.750 83.480 108.830 ;
        RECT 83.950 108.750 84.110 112.730 ;
        RECT 96.030 112.400 96.275 113.350 ;
        RECT 87.160 111.160 87.420 111.480 ;
        RECT 87.210 109.090 87.365 111.160 ;
        RECT 96.030 110.620 96.290 112.400 ;
        RECT 96.030 110.360 96.350 110.620 ;
        RECT 91.770 110.120 92.310 110.230 ;
        RECT 91.770 109.975 97.550 110.120 ;
        RECT 97.710 109.975 97.930 113.960 ;
        RECT 99.965 113.920 100.355 113.960 ;
        RECT 103.315 113.085 103.750 114.420 ;
        RECT 110.725 113.435 110.900 115.280 ;
        RECT 114.590 115.210 115.155 116.800 ;
        RECT 110.725 113.265 115.495 113.435 ;
        RECT 100.890 112.610 101.170 112.645 ;
        RECT 100.470 112.310 101.550 112.610 ;
        RECT 100.890 112.275 101.170 112.310 ;
        RECT 103.325 111.215 103.735 113.085 ;
        RECT 104.955 112.705 105.275 112.965 ;
        RECT 105.040 112.370 105.195 112.705 ;
        RECT 109.965 112.635 110.285 112.895 ;
        RECT 104.970 111.980 105.270 112.370 ;
        RECT 110.050 111.885 110.205 112.635 ;
        RECT 110.480 111.970 110.740 112.290 ;
        RECT 104.400 111.615 104.660 111.695 ;
        RECT 104.400 111.460 106.015 111.615 ;
        RECT 110.000 111.565 110.260 111.885 ;
        RECT 104.400 111.375 104.660 111.460 ;
        RECT 105.860 111.435 106.015 111.460 ;
        RECT 105.860 111.225 106.270 111.435 ;
        RECT 99.200 109.975 99.460 110.010 ;
        RECT 91.770 109.860 99.460 109.975 ;
        RECT 91.770 109.750 92.310 109.860 ;
        RECT 96.805 109.725 99.460 109.860 ;
        RECT 96.805 109.520 97.055 109.725 ;
        RECT 99.200 109.690 99.460 109.725 ;
        RECT 87.125 108.830 87.445 109.090 ;
        RECT 85.665 108.750 86.055 108.825 ;
        RECT 83.220 108.595 86.055 108.750 ;
        RECT 83.220 108.510 83.480 108.595 ;
        RECT 83.950 108.590 84.110 108.595 ;
        RECT 85.665 108.525 86.055 108.595 ;
        RECT 96.770 108.010 97.250 109.520 ;
        RECT 103.345 109.335 103.715 111.215 ;
        RECT 105.950 111.175 106.270 111.225 ;
        RECT 110.525 109.850 110.695 111.970 ;
        RECT 115.325 110.710 115.495 113.265 ;
        RECT 115.250 110.450 115.570 110.710 ;
        RECT 110.450 109.590 110.770 109.850 ;
        RECT 105.400 109.335 105.660 109.360 ;
        RECT 103.345 109.045 105.730 109.335 ;
        RECT 103.345 109.005 103.715 109.045 ;
        RECT 105.400 109.040 105.660 109.045 ;
        RECT 102.935 108.060 103.325 108.135 ;
        RECT 88.890 107.930 89.170 107.965 ;
        RECT 88.560 107.630 89.360 107.930 ;
        RECT 88.890 107.595 89.170 107.630 ;
        RECT 96.740 107.530 97.280 108.010 ;
        RECT 102.805 107.905 103.455 108.060 ;
        RECT 113.790 107.955 114.110 107.975 ;
        RECT 115.820 107.955 116.140 107.975 ;
        RECT 102.935 107.835 103.325 107.905 ;
        RECT 105.740 107.780 106.020 107.815 ;
        RECT 105.730 107.480 106.970 107.780 ;
        RECT 113.790 107.735 116.140 107.955 ;
        RECT 113.790 107.715 114.110 107.735 ;
        RECT 115.820 107.715 116.140 107.735 ;
        RECT 105.740 107.445 106.020 107.480 ;
        RECT 92.840 106.390 97.260 106.870 ;
        RECT 80.135 104.295 80.525 104.335 ;
        RECT 85.730 104.295 85.990 104.345 ;
        RECT 80.135 104.075 85.990 104.295 ;
        RECT 80.135 104.035 80.525 104.075 ;
        RECT 85.730 104.025 85.990 104.075 ;
        RECT 92.840 104.045 93.320 106.390 ;
        RECT 96.675 105.125 96.935 105.210 ;
        RECT 98.855 105.125 99.175 105.175 ;
        RECT 96.675 104.970 99.175 105.125 ;
        RECT 96.675 104.890 96.935 104.970 ;
        RECT 98.855 104.915 99.175 104.970 ;
      LAYER met3 ;
        RECT 113.430 197.890 113.810 198.210 ;
        RECT 116.190 197.890 116.570 198.210 ;
        RECT 113.470 179.215 113.770 197.890 ;
        RECT 116.230 179.845 116.530 197.890 ;
        RECT 116.215 179.515 116.545 179.845 ;
        RECT 113.455 178.885 113.785 179.215 ;
        RECT 85.870 159.620 86.190 160.000 ;
        RECT 85.880 151.565 86.180 159.620 ;
        RECT 85.855 151.215 86.205 151.565 ;
        RECT 80.170 137.750 80.490 138.130 ;
        RECT 1.130 115.450 2.400 116.130 ;
        RECT 13.360 115.450 14.265 115.475 ;
        RECT 1.130 114.595 14.265 115.450 ;
        RECT 1.130 114.000 2.400 114.595 ;
        RECT 13.360 114.570 14.265 114.595 ;
        RECT 51.930 113.205 52.770 113.230 ;
        RECT 13.415 112.415 52.770 113.205 ;
        RECT 51.930 112.390 52.770 112.415 ;
        RECT 80.180 104.360 80.480 137.750 ;
        RECT 100.665 123.755 100.995 124.085 ;
        RECT 91.625 120.860 92.155 120.885 ;
        RECT 91.625 120.380 96.410 120.860 ;
        RECT 91.625 120.355 92.155 120.380 ;
        RECT 93.445 120.070 93.775 120.075 ;
        RECT 93.445 120.060 93.840 120.070 ;
        RECT 93.030 119.760 94.190 120.060 ;
        RECT 93.445 119.750 93.840 119.760 ;
        RECT 93.445 119.745 93.775 119.750 ;
        RECT 95.930 119.270 96.410 120.380 ;
        RECT 100.680 120.180 100.980 123.755 ;
        RECT 104.920 122.210 105.220 122.460 ;
        RECT 104.895 121.860 105.245 122.210 ;
        RECT 98.090 119.880 100.980 120.180 ;
        RECT 98.090 116.925 98.390 119.880 ;
        RECT 98.065 116.575 98.415 116.925 ;
        RECT 98.090 116.370 98.390 116.575 ;
        RECT 100.025 116.280 100.375 116.305 ;
        RECT 103.630 116.280 104.010 116.290 ;
        RECT 99.810 115.980 104.010 116.280 ;
        RECT 99.990 115.955 100.375 115.980 ;
        RECT 103.630 115.970 104.010 115.980 ;
        RECT 95.980 115.715 96.280 115.850 ;
        RECT 95.975 115.410 96.305 115.715 ;
        RECT 99.990 115.660 100.290 115.955 ;
        RECT 104.920 115.680 105.220 121.860 ;
        RECT 106.545 115.680 106.875 115.695 ;
        RECT 93.635 115.380 93.985 115.405 ;
        RECT 94.730 115.380 95.110 115.390 ;
        RECT 95.975 115.385 96.380 115.410 ;
        RECT 93.290 115.080 95.110 115.380 ;
        RECT 95.980 115.110 96.380 115.385 ;
        RECT 104.920 115.380 106.875 115.680 ;
        RECT 106.545 115.365 106.875 115.380 ;
        RECT 93.635 115.055 93.985 115.080 ;
        RECT 94.730 115.070 95.110 115.080 ;
        RECT 96.000 113.665 96.300 115.110 ;
        RECT 97.395 114.605 100.335 114.955 ;
        RECT 95.985 113.335 96.315 113.665 ;
        RECT 85.685 108.825 86.035 108.850 ;
        RECT 85.685 108.525 86.670 108.825 ;
        RECT 85.685 108.500 86.035 108.525 ;
        RECT 86.370 107.930 86.670 108.525 ;
        RECT 88.865 107.930 89.195 107.945 ;
        RECT 86.370 107.630 89.195 107.930 ;
        RECT 88.865 107.615 89.195 107.630 ;
        RECT 80.155 104.010 80.505 104.360 ;
        RECT 93.895 99.355 94.245 99.385 ;
        RECT 97.395 99.355 97.745 114.605 ;
        RECT 99.985 114.220 100.335 114.605 ;
        RECT 99.690 113.920 100.580 114.220 ;
        RECT 99.985 113.895 100.335 113.920 ;
        RECT 100.865 112.610 101.195 112.625 ;
        RECT 100.865 112.310 103.290 112.610 ;
        RECT 104.970 112.350 105.270 112.620 ;
        RECT 100.865 112.295 101.195 112.310 ;
        RECT 102.990 108.160 103.290 112.310 ;
        RECT 104.945 112.000 105.295 112.350 ;
        RECT 102.955 108.135 103.305 108.160 ;
        RECT 102.450 107.835 103.850 108.135 ;
        RECT 102.955 107.810 103.305 107.835 ;
        RECT 104.970 107.780 105.270 112.000 ;
        RECT 105.715 107.780 106.045 107.795 ;
        RECT 104.970 107.480 106.045 107.780 ;
        RECT 105.715 107.465 106.045 107.480 ;
        RECT 93.895 99.005 97.745 99.355 ;
        RECT 93.895 98.975 94.245 99.005 ;
      LAYER met4 ;
        RECT 99.725 220.595 103.490 220.610 ;
        RECT 86.165 220.500 103.490 220.595 ;
        RECT 107.950 220.500 108.250 224.760 ;
        RECT 86.165 220.200 108.250 220.500 ;
        RECT 86.165 220.105 103.490 220.200 ;
        RECT 107.950 220.170 108.250 220.200 ;
        RECT 86.165 173.655 86.655 220.105 ;
        RECT 99.725 220.095 103.490 220.105 ;
        RECT 78.475 173.165 86.655 173.655 ;
        RECT 93.135 215.620 103.865 215.755 ;
        RECT 93.135 215.520 106.660 215.620 ;
        RECT 110.710 215.520 111.010 224.760 ;
        RECT 93.135 215.220 111.010 215.520 ;
        RECT 93.135 215.125 106.660 215.220 ;
        RECT 93.135 214.985 103.865 215.125 ;
        RECT 80.180 138.105 80.480 173.165 ;
        RECT 93.135 168.635 93.905 214.985 ;
        RECT 113.470 198.215 113.770 224.760 ;
        RECT 116.230 198.215 116.530 224.760 ;
        RECT 113.455 197.885 113.785 198.215 ;
        RECT 116.215 197.885 116.545 198.215 ;
        RECT 83.775 167.865 93.905 168.635 ;
        RECT 85.880 159.975 86.180 167.865 ;
        RECT 85.865 159.645 86.195 159.975 ;
        RECT 80.165 137.775 80.495 138.105 ;
        RECT 93.500 120.390 95.810 120.690 ;
        RECT 93.500 120.075 93.800 120.390 ;
        RECT 93.485 119.745 93.815 120.075 ;
        RECT 94.755 115.380 95.085 115.395 ;
        RECT 95.510 115.380 95.810 120.390 ;
        RECT 103.655 115.965 103.985 116.295 ;
        RECT 94.420 115.080 95.810 115.380 ;
        RECT 94.755 115.065 95.085 115.080 ;
        RECT 13.440 113.205 14.240 113.210 ;
        RECT 6.000 112.415 14.240 113.205 ;
        RECT 13.440 112.410 14.240 112.415 ;
        RECT 93.890 99.000 94.250 99.360 ;
        RECT 103.670 99.150 103.970 115.965 ;
        RECT 93.895 93.450 94.245 99.000 ;
        RECT 103.670 98.850 105.340 99.150 ;
        RECT 105.040 95.400 105.340 98.850 ;
        RECT 93.470 53.190 94.370 93.450 ;
        RECT 104.510 70.070 105.410 95.400 ;
        RECT 104.510 69.170 152.710 70.070 ;
        RECT 93.470 52.290 133.390 53.190 ;
        RECT 132.490 1.000 133.390 52.290 ;
        RECT 151.810 1.000 152.710 69.170 ;
  END
END tt_um_analog_example
END LIBRARY

