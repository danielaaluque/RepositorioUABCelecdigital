VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_relax
  CLASS BLOCK ;
  FOREIGN tt_um_relax ;
  ORIGIN 24.865 16.100 ;
  SIZE 37.740 BY 22.930 ;
  PIN ENABLE
    ANTENNAGATEAREA 1.980000 ;
    PORT
      LAYER li1 ;
        RECT -12.300 -14.705 -9.445 -14.485 ;
      LAYER met1 ;
        RECT -11.625 -14.485 -11.345 -14.455 ;
        RECT -14.100 -14.705 -11.000 -14.485 ;
        RECT -11.625 -14.735 -11.345 -14.705 ;
    END
    PORT
      LAYER li1 ;
        RECT -11.980 4.945 -9.125 5.165 ;
      LAYER met1 ;
        RECT -11.750 5.165 -11.470 5.195 ;
        RECT -14.410 4.945 -11.220 5.165 ;
        RECT -11.750 4.915 -11.470 4.945 ;
    END
  END ENABLE
  PIN VGND
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT -12.485 3.975 -2.435 4.885 ;
        RECT -12.340 3.785 -12.170 3.975 ;
        RECT -20.765 -1.265 -8.405 -1.245 ;
        RECT -5.665 -1.265 11.385 -1.255 ;
        RECT -20.765 -1.285 11.385 -1.265 ;
        RECT -20.785 -2.070 11.385 -1.285 ;
        RECT -20.765 -2.155 11.385 -2.070 ;
        RECT -18.020 -2.345 -17.850 -2.155 ;
        RECT -8.810 -2.165 11.385 -2.155 ;
        RECT -8.810 -2.175 -4.940 -2.165 ;
        RECT -8.810 -2.195 -8.665 -2.175 ;
        RECT -8.835 -2.365 -8.665 -2.195 ;
        RECT -2.615 -2.355 -2.445 -2.165 ;
        RECT 6.400 -2.355 6.570 -2.165 ;
        RECT -11.475 -8.845 -4.510 -8.835 ;
        RECT -11.475 -8.855 4.625 -8.845 ;
        RECT -11.475 -8.865 11.585 -8.855 ;
        RECT -20.685 -8.905 11.585 -8.865 ;
        RECT -20.705 -9.690 11.585 -8.905 ;
        RECT -20.685 -9.745 11.585 -9.690 ;
        RECT -20.685 -9.775 -10.285 -9.745 ;
        RECT -8.380 -9.765 -8.235 -9.745 ;
        RECT -4.815 -9.755 11.585 -9.745 ;
        RECT -17.490 -9.965 -17.320 -9.775 ;
        RECT -8.405 -9.935 -8.235 -9.765 ;
        RECT -2.485 -9.945 -2.315 -9.755 ;
        RECT 3.955 -9.765 11.585 -9.755 ;
        RECT 6.600 -9.955 6.770 -9.765 ;
        RECT -12.805 -15.675 -2.535 -14.765 ;
        RECT -12.660 -15.865 -12.490 -15.675 ;
      LAYER li1 ;
        RECT -11.895 3.955 -11.725 4.435 ;
        RECT -11.055 3.955 -10.885 4.435 ;
        RECT -10.215 3.955 -10.045 4.435 ;
        RECT -9.375 3.955 -9.205 4.435 ;
        RECT -12.490 3.785 -5.130 3.955 ;
        RECT -2.795 3.925 -2.505 4.650 ;
        RECT -2.880 3.755 -2.420 3.925 ;
        RECT -20.715 -2.175 -20.425 -1.450 ;
        RECT -17.575 -2.175 -17.405 -1.695 ;
        RECT -16.735 -2.175 -16.565 -1.695 ;
        RECT -15.895 -2.175 -15.725 -1.695 ;
        RECT -15.055 -2.175 -14.885 -1.695 ;
        RECT -20.800 -2.345 -20.340 -2.175 ;
        RECT -18.170 -2.345 -10.810 -2.175 ;
        RECT -8.725 -2.195 -8.470 -1.735 ;
        RECT -7.800 -2.195 -7.630 -1.735 ;
        RECT -6.960 -2.195 -6.790 -1.735 ;
        RECT -6.120 -2.195 -5.950 -1.735 ;
        RECT -5.280 -2.195 -4.975 -1.735 ;
        RECT -2.670 -2.185 -2.395 -1.365 ;
        RECT -1.725 -2.185 -1.555 -1.715 ;
        RECT -0.885 -2.185 -0.715 -1.715 ;
        RECT -0.045 -2.185 0.125 -1.715 ;
        RECT 0.795 -2.185 0.965 -1.715 ;
        RECT 1.635 -2.185 1.805 -1.715 ;
        RECT 2.475 -2.185 2.645 -1.715 ;
        RECT 3.315 -2.185 3.485 -1.715 ;
        RECT 4.155 -2.185 4.445 -1.715 ;
        RECT 6.765 -2.185 7.095 -1.705 ;
        RECT 7.605 -2.185 7.935 -1.705 ;
        RECT 8.445 -2.185 8.775 -1.705 ;
        RECT 9.285 -2.185 9.615 -1.705 ;
        RECT 10.125 -2.185 10.455 -1.705 ;
        RECT 10.965 -2.185 11.295 -1.385 ;
        RECT -8.980 -2.365 -4.840 -2.195 ;
        RECT -2.760 -2.355 4.600 -2.185 ;
        RECT 6.250 -2.355 11.770 -2.185 ;
        RECT -20.635 -9.795 -20.345 -9.070 ;
        RECT -17.045 -9.795 -16.875 -9.315 ;
        RECT -16.205 -9.795 -16.035 -9.315 ;
        RECT -15.365 -9.795 -15.195 -9.315 ;
        RECT -14.525 -9.795 -14.355 -9.315 ;
        RECT -8.295 -9.765 -8.040 -9.305 ;
        RECT -7.370 -9.765 -7.200 -9.305 ;
        RECT -6.530 -9.765 -6.360 -9.305 ;
        RECT -5.690 -9.765 -5.520 -9.305 ;
        RECT -4.850 -9.765 -4.545 -9.305 ;
        RECT -20.720 -9.965 -20.260 -9.795 ;
        RECT -17.640 -9.965 -10.280 -9.795 ;
        RECT -8.550 -9.935 -4.410 -9.765 ;
        RECT -2.540 -9.775 -2.265 -8.955 ;
        RECT -1.595 -9.775 -1.425 -9.305 ;
        RECT -0.755 -9.775 -0.585 -9.305 ;
        RECT 0.085 -9.775 0.255 -9.305 ;
        RECT 0.925 -9.775 1.095 -9.305 ;
        RECT 1.765 -9.775 1.935 -9.305 ;
        RECT 2.605 -9.775 2.775 -9.305 ;
        RECT 3.445 -9.775 3.615 -9.305 ;
        RECT 4.285 -9.775 4.575 -9.305 ;
        RECT -2.630 -9.945 4.730 -9.775 ;
        RECT 6.965 -9.785 7.295 -9.305 ;
        RECT 7.805 -9.785 8.135 -9.305 ;
        RECT 8.645 -9.785 8.975 -9.305 ;
        RECT 9.485 -9.785 9.815 -9.305 ;
        RECT 10.325 -9.785 10.655 -9.305 ;
        RECT 11.165 -9.785 11.495 -8.985 ;
        RECT 6.450 -9.955 11.970 -9.785 ;
        RECT -12.215 -15.695 -12.045 -15.215 ;
        RECT -11.375 -15.695 -11.205 -15.215 ;
        RECT -10.535 -15.695 -10.365 -15.215 ;
        RECT -9.695 -15.695 -9.525 -15.215 ;
        RECT -12.810 -15.865 -5.450 -15.695 ;
        RECT -2.895 -15.705 -2.605 -14.980 ;
        RECT -2.980 -15.875 -2.520 -15.705 ;
      LAYER met1 ;
        RECT -12.490 4.080 -5.130 4.110 ;
        RECT -12.490 3.925 -2.420 4.080 ;
        RECT -21.815 3.785 -21.495 3.840 ;
        RECT -12.490 3.785 -5.130 3.925 ;
        RECT -21.815 3.630 -5.130 3.785 ;
        RECT -21.815 3.580 -21.495 3.630 ;
        RECT -2.880 3.600 -2.420 3.925 ;
        RECT -20.800 -2.040 -10.810 -2.020 ;
        RECT -5.095 -2.040 11.770 -2.030 ;
        RECT -20.800 -2.175 11.770 -2.040 ;
        RECT -23.325 -2.345 -23.065 -2.260 ;
        RECT -20.800 -2.345 -20.340 -2.175 ;
        RECT -23.325 -2.500 -20.340 -2.345 ;
        RECT -18.170 -2.185 11.770 -2.175 ;
        RECT -18.170 -2.195 -4.840 -2.185 ;
        RECT -18.170 -2.500 -10.810 -2.195 ;
        RECT -23.325 -2.580 -23.065 -2.500 ;
        RECT -8.980 -2.520 -4.840 -2.195 ;
        RECT -2.760 -2.510 4.600 -2.185 ;
        RECT 6.250 -2.510 11.770 -2.185 ;
        RECT -10.545 -9.620 -4.410 -9.610 ;
        RECT -10.545 -9.630 4.730 -9.620 ;
        RECT -10.545 -9.640 11.970 -9.630 ;
        RECT -20.720 -9.765 11.970 -9.640 ;
        RECT -20.720 -9.795 -10.280 -9.765 ;
        RECT -22.805 -9.965 -22.545 -9.880 ;
        RECT -20.720 -9.965 -20.260 -9.795 ;
        RECT -22.805 -10.120 -20.260 -9.965 ;
        RECT -17.640 -10.120 -10.280 -9.795 ;
        RECT -8.550 -9.775 11.970 -9.765 ;
        RECT -8.550 -10.090 -4.410 -9.775 ;
        RECT -2.630 -9.785 11.970 -9.775 ;
        RECT -2.630 -10.100 4.730 -9.785 ;
        RECT 6.450 -10.110 11.970 -9.785 ;
        RECT -22.805 -10.200 -22.545 -10.120 ;
        RECT -12.810 -15.550 -2.835 -15.540 ;
        RECT -12.810 -15.695 -2.520 -15.550 ;
        RECT -18.165 -15.865 -17.845 -15.810 ;
        RECT -12.810 -15.865 -5.450 -15.695 ;
        RECT -18.165 -16.020 -5.450 -15.865 ;
        RECT -18.165 -16.070 -17.845 -16.020 ;
        RECT -2.980 -16.030 -2.520 -15.695 ;
      LAYER met2 ;
        RECT -21.785 3.790 -21.525 3.870 ;
        RECT -24.855 3.635 -21.525 3.790 ;
        RECT -24.855 -9.960 -24.700 3.635 ;
        RECT -21.785 3.550 -21.525 3.635 ;
        RECT -23.355 -2.550 -23.035 -2.290 ;
        RECT -23.270 -9.960 -23.115 -2.550 ;
        RECT -22.835 -9.960 -22.515 -9.910 ;
        RECT -24.865 -10.115 -22.515 -9.960 ;
        RECT -24.855 -12.255 -24.700 -10.115 ;
        RECT -23.270 -10.125 -23.115 -10.115 ;
        RECT -22.835 -10.170 -22.515 -10.115 ;
        RECT -24.855 -12.410 -21.225 -12.255 ;
        RECT -24.855 -12.440 -24.700 -12.410 ;
        RECT -21.380 -15.860 -21.225 -12.410 ;
        RECT -18.135 -15.860 -17.875 -15.780 ;
        RECT -21.380 -16.015 -17.875 -15.860 ;
        RECT -18.135 -16.100 -17.875 -16.015 ;
    END
  END VGND
  PIN Q
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER li1 ;
        RECT 8.305 -8.255 8.475 -7.405 ;
        RECT 9.145 -8.255 9.315 -7.405 ;
        RECT 9.985 -8.255 10.155 -7.405 ;
        RECT 10.825 -8.255 10.995 -7.405 ;
        RECT 8.305 -8.425 10.995 -8.255 ;
        RECT 10.740 -8.965 10.995 -8.425 ;
        RECT 8.305 -9.135 10.995 -8.965 ;
        RECT 8.305 -9.615 8.475 -9.135 ;
        RECT 9.145 -9.615 9.315 -9.135 ;
        RECT 9.985 -9.615 10.155 -9.135 ;
        RECT 10.825 -9.615 10.995 -9.135 ;
      LAYER met1 ;
        RECT 10.740 -8.605 10.995 -8.405 ;
        RECT 10.710 -8.635 11.025 -8.605 ;
        RECT 10.535 -8.640 11.205 -8.635 ;
        RECT 10.535 -8.890 12.875 -8.640 ;
        RECT 10.710 -8.895 12.875 -8.890 ;
        RECT 10.710 -8.925 11.025 -8.895 ;
        RECT 10.740 -9.095 10.995 -8.925 ;
    END
  END Q
  PIN Qn
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER li1 ;
        RECT 8.105 -0.655 8.275 0.195 ;
        RECT 8.945 -0.655 9.115 0.195 ;
        RECT 9.785 -0.655 9.955 0.195 ;
        RECT 10.625 -0.655 10.795 0.195 ;
        RECT 8.105 -0.825 10.795 -0.655 ;
        RECT 10.540 -1.365 10.795 -0.825 ;
        RECT 8.105 -1.535 10.795 -1.365 ;
        RECT 8.105 -2.015 8.275 -1.535 ;
        RECT 8.945 -2.015 9.115 -1.535 ;
        RECT 9.785 -2.015 9.955 -1.535 ;
        RECT 10.625 -2.015 10.795 -1.535 ;
      LAYER met1 ;
        RECT 10.510 -1.145 10.825 -1.085 ;
        RECT 10.355 -1.400 12.795 -1.145 ;
        RECT 10.510 -1.465 10.825 -1.400 ;
    END
  END Qn
  PIN C1
    ANTENNAGATEAREA 5.940000 ;
    ANTENNADIFFAREA 5.724000 ;
    PORT
      LAYER li1 ;
        RECT -17.660 -1.185 -14.805 -0.965 ;
        RECT -17.125 -8.215 -16.795 -7.415 ;
        RECT -16.285 -8.215 -15.955 -7.415 ;
        RECT -15.445 -8.215 -15.115 -7.415 ;
        RECT -14.605 -8.215 -14.275 -7.415 ;
        RECT -13.765 -8.215 -13.435 -7.415 ;
        RECT -12.925 -8.215 -12.595 -7.415 ;
        RECT -12.085 -8.215 -11.755 -7.415 ;
        RECT -11.245 -8.215 -10.915 -7.415 ;
        RECT -17.125 -8.415 -10.915 -8.215 ;
        RECT -14.000 -8.805 -13.520 -8.415 ;
        RECT -13.765 -8.975 -13.520 -8.805 ;
        RECT -11.165 -8.975 -10.915 -8.415 ;
        RECT -7.870 -8.775 -5.015 -8.525 ;
        RECT -13.765 -9.225 -10.915 -8.975 ;
        RECT -12.295 -14.115 -11.965 -13.315 ;
        RECT -11.455 -14.115 -11.125 -13.315 ;
        RECT -10.615 -14.115 -10.285 -13.315 ;
        RECT -9.775 -14.115 -9.445 -13.315 ;
        RECT -8.935 -14.115 -8.605 -13.315 ;
        RECT -8.095 -14.115 -7.765 -13.315 ;
        RECT -7.255 -14.115 -6.925 -13.315 ;
        RECT -6.415 -14.115 -6.085 -13.315 ;
        RECT -12.295 -14.315 -6.085 -14.115 ;
        RECT -9.170 -14.705 -8.690 -14.315 ;
        RECT -8.520 -14.705 -6.505 -14.505 ;
        RECT -8.935 -14.875 -8.690 -14.705 ;
        RECT -6.335 -14.875 -6.085 -14.315 ;
        RECT -8.935 -15.125 -6.085 -14.875 ;
      LAYER met1 ;
        RECT -16.290 -0.935 -16.030 -0.915 ;
        RECT -16.565 -0.965 -16.030 -0.935 ;
        RECT -16.850 -1.185 -16.030 -0.965 ;
        RECT -16.565 -1.215 -16.030 -1.185 ;
        RECT -16.290 -1.235 -16.030 -1.215 ;
        RECT -14.030 -8.325 -13.490 -8.295 ;
        RECT -14.350 -8.805 -13.180 -8.325 ;
        RECT -5.970 -8.520 -5.660 -8.495 ;
        RECT -5.980 -8.525 -5.660 -8.520 ;
        RECT -6.405 -8.775 -5.385 -8.525 ;
        RECT -5.980 -8.780 -5.660 -8.775 ;
        RECT -5.970 -8.805 -5.660 -8.780 ;
        RECT -14.030 -8.835 -13.490 -8.805 ;
        RECT -9.200 -14.225 -8.660 -14.195 ;
        RECT -9.450 -14.705 -8.350 -14.225 ;
        RECT -8.140 -14.505 -7.820 -14.475 ;
        RECT -7.420 -14.505 -7.160 -14.475 ;
        RECT -8.140 -14.705 -6.830 -14.505 ;
        RECT -9.200 -14.735 -8.660 -14.705 ;
        RECT -8.140 -14.735 -7.820 -14.705 ;
        RECT -7.420 -14.735 -7.160 -14.705 ;
      LAYER met2 ;
        RECT -16.320 -1.205 -16.000 -0.945 ;
        RECT -16.270 -2.610 -16.050 -1.205 ;
        RECT -16.445 -4.990 -15.870 -2.610 ;
        RECT -16.445 -5.470 -13.520 -4.990 ;
        RECT -16.445 -5.485 -15.870 -5.470 ;
        RECT -14.000 -11.430 -13.520 -5.470 ;
        RECT -9.640 -6.560 -5.950 -6.080 ;
        RECT -9.640 -11.430 -9.160 -6.560 ;
        RECT -5.950 -8.810 -5.690 -8.490 ;
        RECT -5.945 -11.430 -5.695 -8.810 ;
        RECT -14.000 -11.910 -5.690 -11.430 ;
        RECT -9.160 -14.505 -8.680 -11.910 ;
        RECT -8.110 -14.505 -7.850 -14.445 ;
        RECT -9.160 -14.705 -7.850 -14.505 ;
        RECT -9.160 -14.735 -8.680 -14.705 ;
        RECT -8.110 -14.765 -7.850 -14.705 ;
      LAYER met3 ;
        RECT -6.535 -6.080 -6.005 -6.055 ;
        RECT -5.680 -6.080 -5.200 -5.580 ;
        RECT -6.535 -6.560 -5.200 -6.080 ;
        RECT -6.535 -6.585 -6.005 -6.560 ;
        RECT -5.670 -6.570 -5.210 -6.560 ;
    END
  END C1
  PIN C2
    ANTENNAGATEAREA 5.940000 ;
    ANTENNADIFFAREA 5.724000 ;
    PORT
      LAYER li1 ;
        RECT -11.975 5.535 -11.645 6.335 ;
        RECT -11.135 5.535 -10.805 6.335 ;
        RECT -10.295 5.535 -9.965 6.335 ;
        RECT -9.455 5.535 -9.125 6.335 ;
        RECT -8.615 5.535 -8.285 6.335 ;
        RECT -7.775 5.535 -7.445 6.335 ;
        RECT -6.935 5.535 -6.605 6.335 ;
        RECT -6.095 5.535 -5.765 6.335 ;
        RECT -11.975 5.335 -5.765 5.535 ;
        RECT -8.850 4.945 -8.370 5.335 ;
        RECT -8.200 4.945 -6.185 5.145 ;
        RECT -8.615 4.775 -8.370 4.945 ;
        RECT -6.015 4.775 -5.765 5.335 ;
        RECT -8.615 4.525 -5.765 4.775 ;
        RECT -17.655 -0.595 -17.325 0.205 ;
        RECT -16.815 -0.595 -16.485 0.205 ;
        RECT -15.975 -0.595 -15.645 0.205 ;
        RECT -15.135 -0.595 -14.805 0.205 ;
        RECT -14.295 -0.595 -13.965 0.205 ;
        RECT -13.455 -0.595 -13.125 0.205 ;
        RECT -12.615 -0.595 -12.285 0.205 ;
        RECT -11.775 -0.595 -11.445 0.205 ;
        RECT -17.655 -0.795 -11.445 -0.595 ;
        RECT -14.530 -1.185 -14.050 -0.795 ;
        RECT -14.295 -1.355 -14.050 -1.185 ;
        RECT -11.695 -1.355 -11.445 -0.795 ;
        RECT -8.300 -1.205 -5.445 -0.955 ;
        RECT -14.295 -1.605 -11.445 -1.355 ;
        RECT -13.350 -8.805 -11.335 -8.605 ;
      LAYER met1 ;
        RECT -8.850 5.455 -8.370 5.680 ;
        RECT -8.880 4.915 -8.340 5.455 ;
        RECT -7.600 5.145 -7.280 5.175 ;
        RECT -6.665 5.145 -6.405 5.175 ;
        RECT -7.600 4.945 -5.960 5.145 ;
        RECT -7.600 4.915 -7.280 4.945 ;
        RECT -6.665 4.915 -6.405 4.945 ;
        RECT -8.850 4.510 -8.370 4.915 ;
        RECT -14.560 -0.705 -14.020 -0.675 ;
        RECT -14.950 -1.185 -13.560 -0.705 ;
        RECT -7.240 -0.950 -6.930 -0.925 ;
        RECT -7.240 -0.955 -6.920 -0.950 ;
        RECT -14.560 -1.215 -14.020 -1.185 ;
        RECT -7.625 -1.205 -6.745 -0.955 ;
        RECT -7.240 -1.210 -6.920 -1.205 ;
        RECT -7.240 -1.235 -6.930 -1.210 ;
        RECT -12.110 -8.575 -11.850 -8.545 ;
        RECT -12.250 -8.605 -11.850 -8.575 ;
        RECT -12.570 -8.805 -11.650 -8.605 ;
        RECT -12.250 -8.835 -11.850 -8.805 ;
        RECT -12.110 -8.865 -11.850 -8.835 ;
      LAYER met2 ;
        RECT -7.570 5.145 -7.310 5.205 ;
        RECT -8.870 5.020 -7.310 5.145 ;
        RECT -8.880 4.945 -7.310 5.020 ;
        RECT -8.880 4.540 -8.340 4.945 ;
        RECT -7.570 4.885 -7.310 4.945 ;
        RECT -8.850 2.670 -8.370 4.540 ;
        RECT -14.530 2.190 -6.930 2.670 ;
        RECT -14.530 -3.700 -14.050 2.190 ;
        RECT -14.530 -4.180 -11.725 -3.700 ;
        RECT -12.230 -8.955 -11.725 -4.180 ;
        RECT -10.360 -3.720 -9.880 2.190 ;
        RECT -7.205 -0.920 -6.955 2.190 ;
        RECT -7.210 -1.240 -6.950 -0.920 ;
        RECT -10.360 -4.200 -5.155 -3.720 ;
      LAYER met3 ;
        RECT -5.705 -4.225 -5.175 -3.695 ;
        RECT -5.680 -4.820 -5.200 -4.225 ;
    END
  END C2
  OBS
      LAYER nwell ;
        RECT -12.680 6.750 -2.750 6.780 ;
        RECT -12.680 5.175 -2.230 6.750 ;
        RECT -3.070 5.145 -2.230 5.175 ;
        RECT -20.990 0.630 -10.620 0.650 ;
        RECT -5.540 0.630 11.960 0.640 ;
        RECT -20.990 -0.955 11.960 0.630 ;
        RECT -11.510 -0.965 11.960 -0.955 ;
        RECT -11.510 -0.975 -4.650 -0.965 ;
        RECT -10.920 -6.950 -4.220 -6.940 ;
        RECT -10.920 -6.960 4.920 -6.950 ;
        RECT -10.920 -6.970 12.160 -6.960 ;
        RECT -20.910 -8.545 12.160 -6.970 ;
        RECT -20.910 -8.575 -10.090 -8.545 ;
        RECT -4.970 -8.555 12.160 -8.545 ;
        RECT 3.870 -8.565 12.160 -8.555 ;
        RECT -13.000 -12.880 -2.750 -12.870 ;
        RECT -13.000 -14.475 -2.330 -12.880 ;
        RECT -3.170 -14.485 -2.330 -14.475 ;
      LAYER li1 ;
        RECT -12.490 6.505 -5.130 6.675 ;
        RECT -12.400 5.365 -12.145 6.505 ;
        RECT -11.475 5.705 -11.305 6.505 ;
        RECT -10.635 5.705 -10.465 6.505 ;
        RECT -9.795 5.705 -9.625 6.505 ;
        RECT -8.955 5.705 -8.785 6.505 ;
        RECT -8.115 5.705 -7.945 6.505 ;
        RECT -7.275 5.705 -7.105 6.505 ;
        RECT -6.435 5.705 -6.265 6.505 ;
        RECT -5.575 5.365 -5.220 6.505 ;
        RECT -2.880 6.475 -2.420 6.645 ;
        RECT -2.795 5.310 -2.505 6.475 ;
        RECT -12.400 4.605 -8.785 4.775 ;
        RECT -12.400 4.125 -12.065 4.605 ;
        RECT -11.555 4.125 -11.225 4.605 ;
        RECT -10.715 4.125 -10.385 4.605 ;
        RECT -9.875 4.125 -9.545 4.605 ;
        RECT -9.035 4.355 -8.785 4.605 ;
        RECT -5.595 4.355 -5.220 4.775 ;
        RECT -9.035 4.125 -5.220 4.355 ;
        RECT -20.800 0.375 -20.340 0.545 ;
        RECT -18.170 0.375 -10.810 0.545 ;
        RECT -20.715 -0.790 -20.425 0.375 ;
        RECT -18.080 -0.765 -17.825 0.375 ;
        RECT -17.155 -0.425 -16.985 0.375 ;
        RECT -16.315 -0.425 -16.145 0.375 ;
        RECT -15.475 -0.425 -15.305 0.375 ;
        RECT -14.635 -0.425 -14.465 0.375 ;
        RECT -13.795 -0.425 -13.625 0.375 ;
        RECT -12.955 -0.425 -12.785 0.375 ;
        RECT -12.115 -0.425 -11.945 0.375 ;
        RECT -11.255 -0.765 -10.900 0.375 ;
        RECT -8.980 0.355 -4.840 0.525 ;
        RECT -2.760 0.365 4.600 0.535 ;
        RECT 6.250 0.365 11.770 0.535 ;
        RECT -8.725 -0.445 -8.470 0.355 ;
        RECT -8.300 -0.615 -7.970 0.185 ;
        RECT -7.800 -0.445 -7.630 0.355 ;
        RECT -7.460 -0.615 -7.130 0.185 ;
        RECT -6.960 -0.445 -6.790 0.355 ;
        RECT -6.620 -0.615 -6.290 0.185 ;
        RECT -6.120 -0.445 -5.950 0.355 ;
        RECT -5.780 -0.615 -5.450 0.185 ;
        RECT -5.280 -0.445 -4.980 0.355 ;
        RECT -2.670 -0.605 -2.355 0.195 ;
        RECT -2.185 -0.435 -1.935 0.365 ;
        RECT -1.765 -0.605 -1.515 0.195 ;
        RECT -1.345 -0.435 -1.095 0.365 ;
        RECT -0.925 -0.605 -0.675 0.195 ;
        RECT -0.505 -0.435 -0.255 0.365 ;
        RECT -0.085 -0.605 0.165 0.195 ;
        RECT 0.335 -0.435 0.585 0.365 ;
        RECT 0.755 0.025 4.365 0.195 ;
        RECT 0.755 -0.605 1.005 0.025 ;
        RECT -8.895 -0.785 -4.925 -0.615 ;
        RECT -13.880 -1.185 -11.865 -0.985 ;
        RECT -18.080 -1.525 -14.465 -1.355 ;
        RECT -18.080 -2.005 -17.745 -1.525 ;
        RECT -17.235 -2.005 -16.905 -1.525 ;
        RECT -16.395 -2.005 -16.065 -1.525 ;
        RECT -15.555 -2.005 -15.225 -1.525 ;
        RECT -14.715 -1.775 -14.465 -1.525 ;
        RECT -11.275 -1.775 -10.900 -1.355 ;
        RECT -8.895 -1.375 -8.550 -0.785 ;
        RECT -5.245 -1.375 -4.925 -0.785 ;
        RECT -2.670 -0.815 1.005 -0.605 ;
        RECT 1.175 -0.655 1.425 -0.145 ;
        RECT 1.595 -0.485 1.845 0.025 ;
        RECT 2.015 -0.655 2.265 -0.145 ;
        RECT 2.435 -0.485 2.685 0.025 ;
        RECT 2.855 -0.655 3.105 -0.145 ;
        RECT 3.275 -0.485 3.525 0.025 ;
        RECT 3.695 -0.655 3.945 -0.145 ;
        RECT 4.115 -0.485 4.365 0.025 ;
        RECT 6.345 -0.655 6.675 0.195 ;
        RECT 6.845 -0.435 7.015 0.365 ;
        RECT 7.185 -0.655 7.515 0.195 ;
        RECT 7.685 -0.435 7.855 0.365 ;
        RECT 8.445 -0.435 8.775 0.365 ;
        RECT 9.285 -0.435 9.615 0.365 ;
        RECT 10.125 -0.435 10.455 0.365 ;
        RECT 1.175 -0.825 4.515 -0.655 ;
        RECT 6.345 -0.825 7.845 -0.655 ;
        RECT 10.965 -0.785 11.295 0.365 ;
        RECT 3.950 -0.995 4.515 -0.825 ;
        RECT -2.400 -1.195 0.770 -0.995 ;
        RECT 1.040 -1.195 3.780 -0.995 ;
        RECT 3.950 -1.165 4.525 -0.995 ;
        RECT 3.950 -1.365 4.515 -1.165 ;
        RECT 6.390 -1.195 7.490 -0.995 ;
        RECT 7.670 -1.025 7.845 -0.825 ;
        RECT 7.670 -1.195 10.295 -1.025 ;
        RECT 7.670 -1.365 7.845 -1.195 ;
        RECT -8.895 -1.565 -4.925 -1.375 ;
        RECT -2.225 -1.545 4.515 -1.365 ;
        RECT 6.425 -1.535 7.845 -1.365 ;
        RECT -14.715 -2.005 -10.900 -1.775 ;
        RECT -8.300 -2.025 -7.970 -1.565 ;
        RECT -7.460 -2.025 -7.130 -1.565 ;
        RECT -6.620 -2.025 -6.290 -1.565 ;
        RECT -5.780 -2.025 -5.450 -1.565 ;
        RECT -2.225 -2.015 -1.895 -1.545 ;
        RECT -1.385 -2.015 -1.055 -1.545 ;
        RECT -0.545 -2.015 -0.215 -1.545 ;
        RECT 0.295 -2.015 0.625 -1.545 ;
        RECT 1.135 -2.015 1.465 -1.545 ;
        RECT 1.975 -2.015 2.305 -1.545 ;
        RECT 2.815 -2.015 3.145 -1.545 ;
        RECT 3.655 -2.015 3.985 -1.545 ;
        RECT 6.425 -2.015 6.595 -1.535 ;
        RECT 7.265 -2.010 7.435 -1.535 ;
        RECT -20.720 -7.245 -20.260 -7.075 ;
        RECT -17.640 -7.245 -10.280 -7.075 ;
        RECT -8.550 -7.215 -4.410 -7.045 ;
        RECT -20.635 -8.410 -20.345 -7.245 ;
        RECT -17.550 -8.385 -17.295 -7.245 ;
        RECT -16.625 -8.045 -16.455 -7.245 ;
        RECT -15.785 -8.045 -15.615 -7.245 ;
        RECT -14.945 -8.045 -14.775 -7.245 ;
        RECT -14.105 -8.045 -13.935 -7.245 ;
        RECT -13.265 -8.045 -13.095 -7.245 ;
        RECT -12.425 -8.045 -12.255 -7.245 ;
        RECT -11.585 -8.045 -11.415 -7.245 ;
        RECT -10.725 -8.385 -10.370 -7.245 ;
        RECT -8.295 -8.015 -8.040 -7.215 ;
        RECT -7.870 -8.185 -7.540 -7.385 ;
        RECT -7.370 -8.015 -7.200 -7.215 ;
        RECT -7.030 -8.185 -6.700 -7.385 ;
        RECT -6.530 -8.015 -6.360 -7.215 ;
        RECT -6.190 -8.185 -5.860 -7.385 ;
        RECT -5.690 -8.015 -5.520 -7.215 ;
        RECT -5.350 -8.185 -5.020 -7.385 ;
        RECT -4.850 -8.015 -4.550 -7.215 ;
        RECT -2.630 -7.225 4.730 -7.055 ;
        RECT -8.465 -8.355 -4.495 -8.185 ;
        RECT -17.130 -8.805 -14.275 -8.585 ;
        RECT -8.465 -8.945 -8.120 -8.355 ;
        RECT -4.815 -8.945 -4.495 -8.355 ;
        RECT -2.540 -8.195 -2.225 -7.395 ;
        RECT -2.055 -8.025 -1.805 -7.225 ;
        RECT -1.635 -8.195 -1.385 -7.395 ;
        RECT -1.215 -8.025 -0.965 -7.225 ;
        RECT -0.795 -8.195 -0.545 -7.395 ;
        RECT -0.375 -8.025 -0.125 -7.225 ;
        RECT 0.045 -8.195 0.295 -7.395 ;
        RECT 0.465 -8.025 0.715 -7.225 ;
        RECT 6.450 -7.235 11.970 -7.065 ;
        RECT 0.885 -7.565 4.495 -7.395 ;
        RECT 0.885 -8.195 1.135 -7.565 ;
        RECT -2.540 -8.405 1.135 -8.195 ;
        RECT 1.305 -8.245 1.555 -7.735 ;
        RECT 1.725 -8.075 1.975 -7.565 ;
        RECT 2.145 -8.245 2.395 -7.735 ;
        RECT 2.565 -8.075 2.815 -7.565 ;
        RECT 2.985 -8.245 3.235 -7.735 ;
        RECT 3.405 -8.075 3.655 -7.565 ;
        RECT 3.825 -8.245 4.075 -7.735 ;
        RECT 4.245 -8.075 4.495 -7.565 ;
        RECT 1.305 -8.415 4.645 -8.245 ;
        RECT -2.270 -8.785 0.900 -8.585 ;
        RECT 1.170 -8.785 3.910 -8.585 ;
        RECT -17.550 -9.145 -13.935 -8.975 ;
        RECT -17.550 -9.625 -17.215 -9.145 ;
        RECT -16.705 -9.625 -16.375 -9.145 ;
        RECT -15.865 -9.625 -15.535 -9.145 ;
        RECT -15.025 -9.625 -14.695 -9.145 ;
        RECT -14.185 -9.395 -13.935 -9.145 ;
        RECT -10.745 -9.395 -10.370 -8.975 ;
        RECT -8.465 -9.135 -4.495 -8.945 ;
        RECT 4.080 -8.955 4.645 -8.415 ;
        RECT 6.545 -8.255 6.875 -7.405 ;
        RECT 7.045 -8.035 7.215 -7.235 ;
        RECT 7.385 -8.255 7.715 -7.405 ;
        RECT 7.885 -8.035 8.055 -7.235 ;
        RECT 8.645 -8.035 8.975 -7.235 ;
        RECT 9.485 -8.035 9.815 -7.235 ;
        RECT 10.325 -8.035 10.655 -7.235 ;
        RECT 6.545 -8.425 8.045 -8.255 ;
        RECT 11.165 -8.385 11.495 -7.235 ;
        RECT 6.590 -8.795 7.690 -8.595 ;
        RECT 7.870 -8.625 8.045 -8.425 ;
        RECT 7.870 -8.795 10.495 -8.625 ;
        RECT -2.095 -9.135 4.645 -8.955 ;
        RECT 7.870 -8.965 8.045 -8.795 ;
        RECT 6.625 -9.135 8.045 -8.965 ;
        RECT -14.185 -9.625 -10.370 -9.395 ;
        RECT -7.870 -9.595 -7.540 -9.135 ;
        RECT -7.030 -9.595 -6.700 -9.135 ;
        RECT -6.190 -9.595 -5.860 -9.135 ;
        RECT -5.350 -9.595 -5.020 -9.135 ;
        RECT -2.095 -9.605 -1.765 -9.135 ;
        RECT -1.255 -9.605 -0.925 -9.135 ;
        RECT -0.415 -9.605 -0.085 -9.135 ;
        RECT 0.425 -9.605 0.755 -9.135 ;
        RECT 1.265 -9.605 1.595 -9.135 ;
        RECT 2.105 -9.605 2.435 -9.135 ;
        RECT 2.945 -9.605 3.275 -9.135 ;
        RECT 3.785 -9.605 4.115 -9.135 ;
        RECT 6.625 -9.615 6.795 -9.135 ;
        RECT 7.465 -9.610 7.635 -9.135 ;
        RECT -12.810 -13.145 -5.450 -12.975 ;
        RECT -12.720 -14.285 -12.465 -13.145 ;
        RECT -11.795 -13.945 -11.625 -13.145 ;
        RECT -10.955 -13.945 -10.785 -13.145 ;
        RECT -10.115 -13.945 -9.945 -13.145 ;
        RECT -9.275 -13.945 -9.105 -13.145 ;
        RECT -8.435 -13.945 -8.265 -13.145 ;
        RECT -7.595 -13.945 -7.425 -13.145 ;
        RECT -6.755 -13.945 -6.585 -13.145 ;
        RECT -5.895 -14.285 -5.540 -13.145 ;
        RECT -2.980 -13.155 -2.520 -12.985 ;
        RECT -2.895 -14.320 -2.605 -13.155 ;
        RECT -12.720 -15.045 -9.105 -14.875 ;
        RECT -12.720 -15.525 -12.385 -15.045 ;
        RECT -11.875 -15.525 -11.545 -15.045 ;
        RECT -11.035 -15.525 -10.705 -15.045 ;
        RECT -10.195 -15.525 -9.865 -15.045 ;
        RECT -9.355 -15.295 -9.105 -15.045 ;
        RECT -5.915 -15.295 -5.540 -14.875 ;
        RECT -9.355 -15.525 -5.540 -15.295 ;
      LAYER met1 ;
        RECT -23.280 6.800 -2.535 6.830 ;
        RECT -23.280 6.675 -2.420 6.800 ;
        RECT -23.265 0.700 -23.110 6.675 ;
        RECT -12.490 6.350 -5.130 6.675 ;
        RECT -2.880 6.320 -2.420 6.675 ;
        RECT -23.280 0.680 -10.810 0.700 ;
        RECT -5.075 0.680 11.770 0.690 ;
        RECT -23.280 0.545 11.770 0.680 ;
        RECT -21.895 -0.550 -21.740 0.545 ;
        RECT -20.800 0.220 -20.340 0.545 ;
        RECT -18.170 0.535 11.770 0.545 ;
        RECT -18.170 0.525 -4.840 0.535 ;
        RECT -18.170 0.220 -10.810 0.525 ;
        RECT -8.980 0.200 -4.840 0.525 ;
        RECT -2.760 0.210 4.600 0.535 ;
        RECT 6.250 0.210 11.770 0.535 ;
        RECT -21.980 -0.810 -21.660 -0.550 ;
        RECT -5.275 -0.950 -4.895 -0.920 ;
        RECT -12.820 -0.985 -12.500 -0.955 ;
        RECT -13.130 -1.185 -12.240 -0.985 ;
        RECT -5.360 -1.025 -2.520 -0.950 ;
        RECT -1.765 -1.025 -1.535 -0.995 ;
        RECT 2.610 -1.015 2.870 -0.940 ;
        RECT 4.325 -0.995 4.555 -0.935 ;
        RECT 6.950 -0.995 7.180 -0.965 ;
        RECT -12.820 -1.215 -12.500 -1.185 ;
        RECT -5.360 -1.195 -1.065 -1.025 ;
        RECT 2.315 -1.185 3.155 -1.015 ;
        RECT 4.325 -1.165 7.355 -0.995 ;
        RECT -5.360 -1.270 -2.520 -1.195 ;
        RECT -1.765 -1.225 -1.535 -1.195 ;
        RECT 2.610 -1.260 2.870 -1.185 ;
        RECT 4.325 -1.225 4.555 -1.165 ;
        RECT -5.275 -1.300 -4.895 -1.270 ;
        RECT 5.405 -1.310 5.575 -1.165 ;
        RECT 6.950 -1.195 7.180 -1.165 ;
        RECT 5.360 -1.630 5.620 -1.310 ;
        RECT -21.955 -5.210 -21.695 -4.890 ;
        RECT -21.905 -6.920 -21.750 -5.210 ;
        RECT -10.900 -6.900 -4.410 -6.890 ;
        RECT -10.900 -6.910 6.645 -6.900 ;
        RECT -10.900 -6.920 11.970 -6.910 ;
        RECT -21.905 -7.035 11.970 -6.920 ;
        RECT -21.905 -7.075 -10.280 -7.035 ;
        RECT -21.905 -8.985 -21.750 -7.075 ;
        RECT -20.720 -7.400 -20.260 -7.075 ;
        RECT -17.640 -7.400 -10.280 -7.075 ;
        RECT -8.550 -7.055 11.970 -7.035 ;
        RECT -8.550 -7.370 -4.410 -7.055 ;
        RECT -2.630 -7.380 4.730 -7.055 ;
        RECT 6.450 -7.390 11.970 -7.055 ;
        RECT -3.360 -7.820 -3.100 -7.500 ;
        RECT -4.845 -8.530 -4.465 -8.500 ;
        RECT -18.880 -8.585 -18.580 -8.560 ;
        RECT -16.890 -8.585 -16.610 -8.555 ;
        RECT -18.880 -8.890 -16.020 -8.585 ;
        RECT -4.930 -8.850 -3.760 -8.530 ;
        RECT -3.315 -8.585 -3.145 -7.820 ;
        RECT 5.480 -8.030 5.740 -7.710 ;
        RECT -1.635 -8.585 -1.405 -8.555 ;
        RECT -3.315 -8.755 -1.185 -8.585 ;
        RECT 2.380 -8.615 2.700 -8.570 ;
        RECT -1.635 -8.785 -1.405 -8.755 ;
        RECT 2.205 -8.785 2.855 -8.615 ;
        RECT 4.355 -8.625 4.645 -8.595 ;
        RECT 5.525 -8.625 5.695 -8.030 ;
        RECT 7.150 -8.625 7.380 -8.595 ;
        RECT 2.380 -8.830 2.700 -8.785 ;
        RECT 4.355 -8.795 7.595 -8.625 ;
        RECT 4.355 -8.825 4.645 -8.795 ;
        RECT -4.845 -8.880 -4.465 -8.850 ;
        RECT -4.200 -8.860 -3.940 -8.850 ;
        RECT -18.880 -8.920 -18.580 -8.890 ;
        RECT 5.525 -8.970 5.695 -8.795 ;
        RECT 7.150 -8.825 7.380 -8.795 ;
        RECT -21.955 -9.305 -21.695 -8.985 ;
        RECT 5.480 -9.290 5.740 -8.970 ;
        RECT -16.680 -11.385 -16.420 -11.065 ;
        RECT -16.625 -12.820 -16.470 -11.385 ;
        RECT -16.625 -12.830 -5.450 -12.820 ;
        RECT -16.625 -12.975 -2.520 -12.830 ;
        RECT -12.810 -12.985 -2.520 -12.975 ;
        RECT -12.810 -13.300 -5.450 -12.985 ;
        RECT -2.980 -13.310 -2.520 -12.985 ;
      LAYER met2 ;
        RECT -21.950 -0.840 -21.690 -0.520 ;
        RECT -21.900 -4.920 -21.745 -0.840 ;
        RECT -12.790 -1.245 -12.530 -0.925 ;
        RECT 2.580 -1.230 2.900 -0.970 ;
        RECT -12.760 -3.065 -12.560 -1.245 ;
        RECT -11.980 -3.065 -11.700 -3.030 ;
        RECT -12.760 -3.365 -11.690 -3.065 ;
        RECT -11.980 -3.400 -11.700 -3.365 ;
        RECT -21.985 -5.180 -21.665 -4.920 ;
        RECT 2.655 -6.055 2.825 -1.230 ;
        RECT 5.330 -1.600 5.650 -1.340 ;
        RECT 3.735 -3.130 4.035 -3.020 ;
        RECT 5.405 -3.130 5.575 -1.600 ;
        RECT 3.735 -3.305 5.580 -3.130 ;
        RECT 3.735 -3.410 4.035 -3.305 ;
        RECT 5.405 -4.235 5.575 -3.305 ;
        RECT 5.340 -4.625 5.640 -4.235 ;
        RECT 1.910 -6.230 2.190 -6.195 ;
        RECT 2.655 -6.225 5.695 -6.055 ;
        RECT -3.320 -6.530 2.200 -6.230 ;
        RECT -3.315 -7.530 -3.145 -6.530 ;
        RECT 1.910 -6.565 2.190 -6.530 ;
        RECT -3.390 -7.790 -3.070 -7.530 ;
        RECT 5.525 -7.740 5.695 -6.225 ;
        RECT 5.450 -8.000 5.770 -7.740 ;
        RECT -18.870 -8.590 -18.590 -8.555 ;
        RECT -18.910 -8.890 -18.550 -8.590 ;
        RECT -4.230 -8.615 -3.910 -8.570 ;
        RECT 2.410 -8.615 2.670 -8.540 ;
        RECT -4.230 -8.785 2.670 -8.615 ;
        RECT -4.230 -8.830 -3.910 -8.785 ;
        RECT 2.410 -8.860 2.670 -8.785 ;
        RECT -18.870 -8.925 -18.590 -8.890 ;
        RECT -21.985 -9.275 -21.665 -9.015 ;
        RECT 5.450 -9.260 5.770 -9.000 ;
        RECT -21.900 -11.150 -21.745 -9.275 ;
        RECT -3.595 -10.885 -3.205 -10.820 ;
        RECT 5.525 -10.885 5.695 -9.260 ;
        RECT -3.595 -11.055 5.695 -10.885 ;
        RECT -16.710 -11.150 -16.390 -11.095 ;
        RECT -3.595 -11.120 -3.205 -11.055 ;
        RECT -21.900 -11.305 -16.390 -11.150 ;
        RECT -16.710 -11.355 -16.390 -11.305 ;
      LAYER met3 ;
        RECT -12.005 -3.065 -11.675 -3.050 ;
        RECT 3.710 -3.065 4.060 -3.040 ;
        RECT -12.005 -3.365 4.550 -3.065 ;
        RECT -12.005 -3.380 -11.675 -3.365 ;
        RECT 3.710 -3.390 4.060 -3.365 ;
        RECT 5.315 -4.605 5.665 -4.255 ;
        RECT 1.885 -6.230 2.215 -6.215 ;
        RECT 5.340 -6.230 5.640 -4.605 ;
        RECT 1.885 -6.530 5.640 -6.230 ;
        RECT 1.885 -6.545 2.215 -6.530 ;
        RECT -18.895 -8.905 -18.565 -8.575 ;
        RECT -18.880 -10.820 -18.580 -8.905 ;
        RECT -3.575 -10.820 -3.225 -10.795 ;
        RECT -18.880 -11.120 -3.225 -10.820 ;
        RECT -3.575 -11.145 -3.225 -11.120 ;
  END
END tt_um_relax
END LIBRARY

