VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_relax
  CLASS BLOCK ;
  FOREIGN tt_um_relax ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 146.590 224.760 146.890 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 141.070 224.760 141.370 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 5.940000 ;
    ANTENNADIFFAREA 5.724000 ;
    PORT
      LAYER li1 ;
        RECT 86.885 127.735 87.215 128.535 ;
        RECT 87.725 127.735 88.055 128.535 ;
        RECT 88.565 127.735 88.895 128.535 ;
        RECT 89.405 127.735 89.735 128.535 ;
        RECT 90.245 127.735 90.575 128.535 ;
        RECT 91.085 127.735 91.415 128.535 ;
        RECT 91.925 127.735 92.255 128.535 ;
        RECT 92.765 127.735 93.095 128.535 ;
        RECT 86.885 127.535 93.095 127.735 ;
        RECT 90.010 127.145 90.490 127.535 ;
        RECT 90.660 127.145 92.675 127.345 ;
        RECT 90.245 126.975 90.490 127.145 ;
        RECT 92.845 126.975 93.095 127.535 ;
        RECT 90.245 126.725 93.095 126.975 ;
        RECT 87.545 120.735 87.875 121.535 ;
        RECT 88.385 120.735 88.715 121.535 ;
        RECT 89.225 120.735 89.555 121.535 ;
        RECT 90.065 120.735 90.395 121.535 ;
        RECT 90.905 120.735 91.235 121.535 ;
        RECT 91.745 120.735 92.075 121.535 ;
        RECT 92.585 120.735 92.915 121.535 ;
        RECT 93.425 120.735 93.755 121.535 ;
        RECT 87.545 120.535 93.755 120.735 ;
        RECT 90.670 120.145 91.150 120.535 ;
        RECT 90.905 119.975 91.150 120.145 ;
        RECT 93.505 119.975 93.755 120.535 ;
        RECT 98.200 120.145 101.055 120.395 ;
        RECT 90.905 119.725 93.755 119.975 ;
        RECT 91.320 113.145 93.335 113.345 ;
      LAYER met1 ;
        RECT 90.040 127.480 90.440 127.640 ;
        RECT 90.850 127.480 91.240 127.530 ;
        RECT 90.040 127.350 91.240 127.480 ;
        RECT 90.040 127.320 94.940 127.350 ;
        RECT 90.040 127.240 90.440 127.320 ;
        RECT 90.850 127.145 94.940 127.320 ;
        RECT 90.850 127.080 91.240 127.145 ;
        RECT 94.720 125.970 94.940 127.145 ;
        RECT 102.880 125.970 103.780 126.000 ;
        RECT 94.720 125.070 103.780 125.970 ;
        RECT 94.720 122.750 94.940 125.070 ;
        RECT 102.880 125.040 103.780 125.070 ;
        RECT 94.670 122.490 94.990 122.750 ;
        RECT 94.700 121.040 94.960 121.090 ;
        RECT 90.770 120.820 96.430 121.040 ;
        RECT 90.770 120.590 90.990 120.820 ;
        RECT 94.700 120.770 94.960 120.820 ;
        RECT 90.650 120.130 91.110 120.590 ;
        RECT 96.175 120.400 96.430 120.820 ;
        RECT 98.320 120.400 98.810 120.520 ;
        RECT 96.175 120.145 98.810 120.400 ;
        RECT 96.175 119.885 96.430 120.145 ;
        RECT 98.320 120.050 98.810 120.145 ;
        RECT 96.175 119.565 96.435 119.885 ;
        RECT 92.415 114.010 92.675 114.330 ;
        RECT 92.415 113.460 92.670 114.010 ;
        RECT 92.310 113.010 92.750 113.460 ;
      LAYER met2 ;
        RECT 129.025 125.970 129.875 125.990 ;
        RECT 102.850 125.070 129.900 125.970 ;
        RECT 129.025 125.050 129.875 125.070 ;
        RECT 94.700 122.460 94.960 122.780 ;
        RECT 94.720 121.060 94.940 122.460 ;
        RECT 94.670 120.800 94.990 121.060 ;
        RECT 96.145 119.595 96.465 119.855 ;
        RECT 92.420 115.840 92.675 115.845 ;
        RECT 96.180 115.840 96.435 119.595 ;
        RECT 92.420 115.585 96.435 115.840 ;
        RECT 92.420 114.300 92.675 115.585 ;
        RECT 92.385 114.040 92.705 114.300 ;
      LAYER met3 ;
        RECT 129.000 125.070 141.600 125.970 ;
        RECT 140.700 20.080 141.600 125.070 ;
        RECT 140.700 19.180 152.710 20.080 ;
        RECT 151.810 5.115 152.710 19.180 ;
        RECT 151.785 4.225 152.735 5.115 ;
        RECT 151.810 4.220 152.710 4.225 ;
      LAYER met4 ;
        RECT 151.810 0.000 152.710 5.120 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 5.940000 ;
    ANTENNADIFFAREA 5.724000 ;
    PORT
      LAYER li1 ;
        RECT 87.540 120.145 90.395 120.365 ;
        RECT 87.545 113.735 87.875 114.535 ;
        RECT 88.385 113.735 88.715 114.535 ;
        RECT 89.225 113.735 89.555 114.535 ;
        RECT 90.065 113.735 90.395 114.535 ;
        RECT 90.905 113.735 91.235 114.535 ;
        RECT 91.745 113.735 92.075 114.535 ;
        RECT 92.585 113.735 92.915 114.535 ;
        RECT 93.425 113.735 93.755 114.535 ;
        RECT 87.545 113.535 93.755 113.735 ;
        RECT 90.670 113.145 91.150 113.535 ;
        RECT 90.905 112.975 91.150 113.145 ;
        RECT 93.505 112.975 93.755 113.535 ;
        RECT 98.210 113.145 101.065 113.395 ;
        RECT 90.905 112.725 93.755 112.975 ;
        RECT 86.835 108.245 87.165 109.045 ;
        RECT 87.675 108.245 88.005 109.045 ;
        RECT 88.515 108.245 88.845 109.045 ;
        RECT 89.355 108.245 89.685 109.045 ;
        RECT 90.195 108.245 90.525 109.045 ;
        RECT 91.035 108.245 91.365 109.045 ;
        RECT 91.875 108.245 92.205 109.045 ;
        RECT 92.715 108.245 93.045 109.045 ;
        RECT 86.835 108.045 93.045 108.245 ;
        RECT 89.960 107.655 90.440 108.045 ;
        RECT 90.610 107.655 92.625 107.855 ;
        RECT 90.195 107.485 90.440 107.655 ;
        RECT 92.795 107.485 93.045 108.045 ;
        RECT 90.195 107.235 93.045 107.485 ;
      LAYER met1 ;
        RECT 87.635 119.900 87.885 120.395 ;
        RECT 87.600 119.640 87.920 119.900 ;
        RECT 90.670 113.130 91.140 113.580 ;
        RECT 98.370 113.400 98.800 113.480 ;
        RECT 96.235 113.145 98.800 113.400 ;
        RECT 87.600 112.860 87.920 112.865 ;
        RECT 90.790 112.860 91.040 113.130 ;
        RECT 94.850 112.860 95.170 112.865 ;
        RECT 96.235 112.860 96.490 113.145 ;
        RECT 98.370 113.050 98.800 113.145 ;
        RECT 87.600 112.610 96.495 112.860 ;
        RECT 87.600 112.605 87.920 112.610 ;
        RECT 94.850 112.605 95.170 112.610 ;
        RECT 94.850 110.340 95.170 110.600 ;
        RECT 94.885 109.300 95.135 110.340 ;
        RECT 94.885 108.400 99.960 109.300 ;
        RECT 90.000 107.940 90.370 108.090 ;
        RECT 90.000 107.850 91.640 107.940 ;
        RECT 94.885 107.850 95.135 108.400 ;
        RECT 90.000 107.720 95.135 107.850 ;
        RECT 91.180 107.655 95.135 107.720 ;
        RECT 91.180 107.540 91.640 107.655 ;
      LAYER met2 ;
        RECT 87.630 119.610 87.890 119.930 ;
        RECT 87.635 112.895 87.885 119.610 ;
        RECT 87.630 112.575 87.890 112.895 ;
        RECT 94.880 112.575 95.140 112.895 ;
        RECT 94.885 110.630 95.135 112.575 ;
        RECT 94.880 110.310 95.140 110.630 ;
        RECT 99.030 65.595 99.930 109.330 ;
        RECT 99.010 64.745 99.950 65.595 ;
        RECT 99.030 64.720 99.930 64.745 ;
      LAYER met3 ;
        RECT 99.030 52.030 99.930 65.620 ;
        RECT 99.030 51.130 133.390 52.030 ;
        RECT 132.490 3.835 133.390 51.130 ;
        RECT 132.465 2.945 133.415 3.835 ;
        RECT 132.490 2.940 133.390 2.945 ;
      LAYER met4 ;
        RECT 132.490 0.000 133.390 3.840 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 113.170 0.000 114.070 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 93.850 0.000 94.750 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 74.530 0.000 75.430 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.210 0.000 56.110 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 35.890 0.000 36.790 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 16.570 0.000 17.470 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 138.310 224.760 138.610 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 135.550 224.760 135.850 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 130.030 224.760 130.330 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 127.270 224.760 127.570 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 124.510 224.760 124.810 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.990 224.760 119.290 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER li1 ;
        RECT 116.875 113.685 117.045 114.535 ;
        RECT 117.715 113.685 117.885 114.535 ;
        RECT 118.555 113.685 118.725 114.535 ;
        RECT 119.395 113.685 119.565 114.535 ;
        RECT 116.875 113.515 119.565 113.685 ;
        RECT 119.310 112.975 119.565 113.515 ;
        RECT 116.875 112.805 119.565 112.975 ;
        RECT 116.875 112.325 117.045 112.805 ;
        RECT 117.715 112.325 117.885 112.805 ;
        RECT 118.555 112.325 118.725 112.805 ;
        RECT 119.395 112.325 119.565 112.805 ;
      LAYER met1 ;
        RECT 128.970 137.100 129.330 137.400 ;
        RECT 119.250 113.340 119.610 113.430 ;
        RECT 129.000 113.340 129.300 137.100 ;
        RECT 119.250 113.140 129.300 113.340 ;
        RECT 119.250 113.060 119.610 113.140 ;
      LAYER met2 ;
        RECT 129.010 209.310 129.290 209.345 ;
        RECT 129.000 137.070 129.300 209.310 ;
      LAYER met3 ;
        RECT 116.190 223.010 116.570 223.330 ;
        RECT 116.230 209.310 116.530 223.010 ;
        RECT 128.985 209.310 129.315 209.325 ;
        RECT 116.230 209.010 129.315 209.310 ;
        RECT 128.985 208.995 129.315 209.010 ;
      LAYER met4 ;
        RECT 116.230 223.335 116.530 225.760 ;
        RECT 116.215 223.005 116.545 223.335 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER li1 ;
        RECT 116.885 120.685 117.055 121.535 ;
        RECT 117.725 120.685 117.895 121.535 ;
        RECT 118.565 120.685 118.735 121.535 ;
        RECT 119.405 120.685 119.575 121.535 ;
        RECT 116.885 120.515 119.575 120.685 ;
        RECT 119.320 119.975 119.575 120.515 ;
        RECT 116.885 119.805 119.575 119.975 ;
        RECT 116.885 119.325 117.055 119.805 ;
        RECT 117.725 119.325 117.895 119.805 ;
        RECT 118.565 119.325 118.735 119.805 ;
        RECT 119.405 119.325 119.575 119.805 ;
      LAYER met1 ;
        RECT 126.380 154.940 126.740 155.240 ;
        RECT 119.220 120.330 119.650 120.440 ;
        RECT 126.410 120.330 126.710 154.940 ;
        RECT 119.220 120.100 126.710 120.330 ;
        RECT 119.220 120.010 119.650 120.100 ;
      LAYER met2 ;
        RECT 126.410 204.550 126.710 204.560 ;
        RECT 126.375 204.270 126.745 204.550 ;
        RECT 126.410 154.910 126.710 204.270 ;
      LAYER met3 ;
        RECT 113.430 222.390 113.810 222.710 ;
        RECT 113.470 204.560 113.770 222.390 ;
        RECT 126.395 204.560 126.725 204.575 ;
        RECT 113.470 204.260 126.725 204.560 ;
        RECT 126.395 204.245 126.725 204.260 ;
      LAYER met4 ;
        RECT 113.470 222.715 113.770 225.760 ;
        RECT 113.455 222.385 113.785 222.715 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.980000 ;
    PORT
      LAYER li1 ;
        RECT 86.880 127.145 89.735 127.365 ;
      LAYER met1 ;
        RECT 84.230 133.870 84.490 134.190 ;
        RECT 84.235 126.890 84.485 133.870 ;
        RECT 87.870 127.050 88.300 127.440 ;
        RECT 87.970 126.890 88.220 127.050 ;
        RECT 84.235 126.640 88.220 126.890 ;
      LAYER met2 ;
        RECT 110.710 166.180 111.010 166.190 ;
        RECT 110.675 165.900 111.045 166.180 ;
        RECT 110.710 136.455 111.010 165.900 ;
        RECT 84.235 136.205 111.015 136.455 ;
        RECT 84.235 134.160 84.485 136.205 ;
        RECT 84.200 133.900 84.520 134.160 ;
      LAYER met3 ;
        RECT 110.670 222.450 111.050 222.770 ;
        RECT 110.710 166.205 111.010 222.450 ;
        RECT 110.695 165.875 111.025 166.205 ;
      LAYER met4 ;
        RECT 110.710 222.775 111.010 225.760 ;
        RECT 110.695 222.445 111.025 222.775 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.980000 ;
    PORT
      LAYER li1 ;
        RECT 86.830 107.655 89.685 107.875 ;
      LAYER met1 ;
        RECT 83.985 107.870 84.305 107.895 ;
        RECT 86.990 107.870 87.430 107.950 ;
        RECT 83.985 107.655 87.430 107.870 ;
        RECT 83.985 107.635 84.305 107.655 ;
        RECT 86.990 107.530 87.430 107.655 ;
      LAYER met2 ;
        RECT 81.365 121.055 81.665 121.445 ;
        RECT 81.405 107.875 81.620 121.055 ;
        RECT 84.015 107.875 84.275 107.925 ;
        RECT 81.405 107.660 84.275 107.875 ;
        RECT 84.015 107.605 84.275 107.660 ;
      LAYER met3 ;
        RECT 107.910 222.270 108.290 222.590 ;
        RECT 107.950 158.050 108.250 222.270 ;
        RECT 81.365 157.750 108.250 158.050 ;
        RECT 81.365 121.425 81.665 157.750 ;
        RECT 81.340 121.075 81.690 121.425 ;
      LAYER met4 ;
        RECT 107.950 222.595 108.250 225.760 ;
        RECT 107.935 222.265 108.265 222.595 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 105.190 224.760 105.490 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 102.430 224.760 102.730 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 96.910 224.760 97.210 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 49.990 224.760 50.290 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 47.230 224.760 47.530 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 41.710 224.760 42.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 38.950 224.760 39.250 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 36.190 224.760 36.490 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 30.670 224.760 30.970 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 72.070 224.760 72.370 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 69.310 224.760 69.610 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 63.790 224.760 64.090 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 61.030 224.760 61.330 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 58.270 224.760 58.570 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 52.750 224.760 53.050 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 94.150 224.760 94.450 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 91.390 224.760 91.690 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 85.870 224.760 86.170 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 83.110 224.760 83.410 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 80.350 224.760 80.650 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 74.830 224.760 75.130 225.760 ;
    END
  END uo_out[7]
  PIN VDPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 85.340 127.375 93.920 128.980 ;
        RECT 84.360 120.375 120.740 121.980 ;
        RECT 84.340 113.375 120.730 114.980 ;
        RECT 85.330 107.885 93.870 109.490 ;
      LAYER li1 ;
        RECT 85.530 128.705 85.990 128.875 ;
        RECT 86.370 128.705 93.730 128.875 ;
        RECT 85.615 127.540 85.905 128.705 ;
        RECT 86.460 127.565 86.715 128.705 ;
        RECT 87.385 127.905 87.555 128.705 ;
        RECT 88.225 127.905 88.395 128.705 ;
        RECT 89.065 127.905 89.235 128.705 ;
        RECT 89.905 127.905 90.075 128.705 ;
        RECT 90.745 127.905 90.915 128.705 ;
        RECT 91.585 127.905 91.755 128.705 ;
        RECT 92.425 127.905 92.595 128.705 ;
        RECT 93.285 127.565 93.640 128.705 ;
        RECT 84.550 121.705 85.010 121.875 ;
        RECT 87.030 121.705 94.390 121.875 ;
        RECT 97.520 121.705 101.660 121.875 ;
        RECT 104.540 121.705 111.900 121.875 ;
        RECT 115.030 121.705 120.550 121.875 ;
        RECT 84.635 120.540 84.925 121.705 ;
        RECT 87.120 120.565 87.375 121.705 ;
        RECT 88.045 120.905 88.215 121.705 ;
        RECT 88.885 120.905 89.055 121.705 ;
        RECT 89.725 120.905 89.895 121.705 ;
        RECT 90.565 120.905 90.735 121.705 ;
        RECT 91.405 120.905 91.575 121.705 ;
        RECT 92.245 120.905 92.415 121.705 ;
        RECT 93.085 120.905 93.255 121.705 ;
        RECT 93.945 120.565 94.300 121.705 ;
        RECT 97.775 120.905 98.030 121.705 ;
        RECT 98.700 120.905 98.870 121.705 ;
        RECT 99.540 120.905 99.710 121.705 ;
        RECT 100.380 120.905 100.550 121.705 ;
        RECT 101.220 120.905 101.520 121.705 ;
        RECT 105.115 120.905 105.365 121.705 ;
        RECT 105.955 120.905 106.205 121.705 ;
        RECT 106.795 120.905 107.045 121.705 ;
        RECT 107.635 120.905 107.885 121.705 ;
        RECT 115.625 120.905 115.795 121.705 ;
        RECT 116.465 120.905 116.635 121.705 ;
        RECT 117.225 120.905 117.555 121.705 ;
        RECT 118.065 120.905 118.395 121.705 ;
        RECT 118.905 120.905 119.235 121.705 ;
        RECT 119.745 120.555 120.075 121.705 ;
        RECT 84.530 114.705 84.990 114.875 ;
        RECT 87.030 114.705 94.390 114.875 ;
        RECT 97.530 114.705 101.670 114.875 ;
        RECT 104.530 114.705 111.890 114.875 ;
        RECT 115.020 114.705 120.540 114.875 ;
        RECT 84.615 113.540 84.905 114.705 ;
        RECT 87.120 113.565 87.375 114.705 ;
        RECT 88.045 113.905 88.215 114.705 ;
        RECT 88.885 113.905 89.055 114.705 ;
        RECT 89.725 113.905 89.895 114.705 ;
        RECT 90.565 113.905 90.735 114.705 ;
        RECT 91.405 113.905 91.575 114.705 ;
        RECT 92.245 113.905 92.415 114.705 ;
        RECT 93.085 113.905 93.255 114.705 ;
        RECT 93.945 113.565 94.300 114.705 ;
        RECT 97.785 113.905 98.040 114.705 ;
        RECT 98.710 113.905 98.880 114.705 ;
        RECT 99.550 113.905 99.720 114.705 ;
        RECT 100.390 113.905 100.560 114.705 ;
        RECT 101.230 113.905 101.530 114.705 ;
        RECT 105.105 113.905 105.355 114.705 ;
        RECT 105.945 113.905 106.195 114.705 ;
        RECT 106.785 113.905 107.035 114.705 ;
        RECT 107.625 113.905 107.875 114.705 ;
        RECT 115.615 113.905 115.785 114.705 ;
        RECT 116.455 113.905 116.625 114.705 ;
        RECT 117.215 113.905 117.545 114.705 ;
        RECT 118.055 113.905 118.385 114.705 ;
        RECT 118.895 113.905 119.225 114.705 ;
        RECT 119.735 113.555 120.065 114.705 ;
        RECT 85.520 109.215 85.980 109.385 ;
        RECT 86.320 109.215 93.680 109.385 ;
        RECT 85.605 108.050 85.895 109.215 ;
        RECT 86.410 108.075 86.665 109.215 ;
        RECT 87.335 108.415 87.505 109.215 ;
        RECT 88.175 108.415 88.345 109.215 ;
        RECT 89.015 108.415 89.185 109.215 ;
        RECT 89.855 108.415 90.025 109.215 ;
        RECT 90.695 108.415 90.865 109.215 ;
        RECT 91.535 108.415 91.705 109.215 ;
        RECT 92.375 108.415 92.545 109.215 ;
        RECT 93.235 108.075 93.590 109.215 ;
      LAYER met1 ;
        RECT 85.530 128.930 93.730 129.030 ;
        RECT 85.520 128.550 93.730 128.930 ;
        RECT 85.520 127.950 86.000 128.550 ;
        RECT 85.490 127.470 86.030 127.950 ;
        RECT 85.520 123.760 86.000 124.990 ;
        RECT 84.110 123.280 86.000 123.760 ;
        RECT 85.520 122.030 86.000 123.280 ;
        RECT 84.550 121.550 120.550 122.030 ;
        RECT 85.520 120.720 86.000 121.550 ;
        RECT 85.490 120.240 86.030 120.720 ;
        RECT 85.520 115.030 86.000 117.870 ;
        RECT 84.530 114.555 120.540 115.030 ;
        RECT 84.530 114.550 84.990 114.555 ;
        RECT 85.520 113.380 86.000 114.555 ;
        RECT 87.030 114.550 94.390 114.555 ;
        RECT 97.530 114.550 101.670 114.555 ;
        RECT 104.530 114.550 111.890 114.555 ;
        RECT 115.020 114.550 120.540 114.555 ;
        RECT 85.490 112.900 86.030 113.380 ;
        RECT 85.520 109.540 86.000 110.780 ;
        RECT 85.520 109.060 93.680 109.540 ;
      LAYER met2 ;
        RECT 85.520 124.960 86.000 127.980 ;
        RECT 85.490 124.480 86.030 124.960 ;
        RECT 45.440 124.020 57.260 124.060 ;
        RECT 45.440 123.885 70.320 124.020 ;
        RECT 45.440 123.760 78.475 123.885 ;
        RECT 84.140 123.760 84.620 123.790 ;
        RECT 45.440 123.280 84.620 123.760 ;
        RECT 45.440 123.155 78.475 123.280 ;
        RECT 84.140 123.250 84.620 123.280 ;
        RECT 45.440 123.020 70.320 123.155 ;
        RECT 45.440 122.985 57.260 123.020 ;
        RECT 85.520 117.840 86.000 120.750 ;
        RECT 85.490 117.360 86.030 117.840 ;
        RECT 85.520 110.750 86.000 113.410 ;
        RECT 85.490 110.270 86.030 110.750 ;
      LAYER met3 ;
        RECT 45.460 124.060 46.585 124.085 ;
        RECT 1.225 122.985 46.585 124.060 ;
        RECT 45.460 122.960 46.585 122.985 ;
      LAYER met4 ;
        RECT 1.000 5.000 3.000 220.760 ;
    END
  END VDPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 85.535 126.175 93.725 127.085 ;
        RECT 86.520 125.985 86.690 126.175 ;
        RECT 84.545 119.175 120.165 120.085 ;
        RECT 87.180 118.985 87.350 119.175 ;
        RECT 97.690 119.155 97.835 119.175 ;
        RECT 97.665 118.985 97.835 119.155 ;
        RECT 104.685 118.985 104.855 119.175 ;
        RECT 115.180 118.985 115.350 119.175 ;
        RECT 84.545 112.175 120.155 113.085 ;
        RECT 87.180 111.985 87.350 112.175 ;
        RECT 97.700 112.155 97.845 112.175 ;
        RECT 97.675 111.985 97.845 112.155 ;
        RECT 104.675 111.985 104.845 112.175 ;
        RECT 115.170 111.985 115.340 112.175 ;
        RECT 85.545 107.555 93.675 107.595 ;
        RECT 85.535 106.770 93.675 107.555 ;
        RECT 85.545 106.685 93.675 106.770 ;
        RECT 86.470 106.495 86.640 106.685 ;
      LAYER li1 ;
        RECT 85.615 126.155 85.905 126.880 ;
        RECT 86.965 126.155 87.135 126.635 ;
        RECT 87.805 126.155 87.975 126.635 ;
        RECT 88.645 126.155 88.815 126.635 ;
        RECT 89.485 126.155 89.655 126.635 ;
        RECT 85.530 125.985 85.990 126.155 ;
        RECT 86.370 125.985 93.730 126.155 ;
        RECT 84.635 119.155 84.925 119.880 ;
        RECT 87.625 119.155 87.795 119.635 ;
        RECT 88.465 119.155 88.635 119.635 ;
        RECT 89.305 119.155 89.475 119.635 ;
        RECT 90.145 119.155 90.315 119.635 ;
        RECT 97.775 119.155 98.030 119.615 ;
        RECT 98.700 119.155 98.870 119.615 ;
        RECT 99.540 119.155 99.710 119.615 ;
        RECT 100.380 119.155 100.550 119.615 ;
        RECT 101.220 119.155 101.525 119.615 ;
        RECT 104.630 119.155 104.905 119.975 ;
        RECT 105.575 119.155 105.745 119.625 ;
        RECT 106.415 119.155 106.585 119.625 ;
        RECT 107.255 119.155 107.425 119.625 ;
        RECT 108.095 119.155 108.265 119.625 ;
        RECT 108.935 119.155 109.105 119.625 ;
        RECT 109.775 119.155 109.945 119.625 ;
        RECT 110.615 119.155 110.785 119.625 ;
        RECT 111.455 119.155 111.745 119.625 ;
        RECT 115.545 119.155 115.875 119.635 ;
        RECT 116.385 119.155 116.715 119.635 ;
        RECT 117.225 119.155 117.555 119.635 ;
        RECT 118.065 119.155 118.395 119.635 ;
        RECT 118.905 119.155 119.235 119.635 ;
        RECT 119.745 119.155 120.075 119.955 ;
        RECT 84.550 118.985 85.010 119.155 ;
        RECT 87.030 118.985 94.390 119.155 ;
        RECT 97.520 118.985 101.660 119.155 ;
        RECT 104.540 118.985 111.900 119.155 ;
        RECT 115.030 118.985 120.550 119.155 ;
        RECT 84.615 112.155 84.905 112.880 ;
        RECT 87.625 112.155 87.795 112.635 ;
        RECT 88.465 112.155 88.635 112.635 ;
        RECT 89.305 112.155 89.475 112.635 ;
        RECT 90.145 112.155 90.315 112.635 ;
        RECT 97.785 112.155 98.040 112.615 ;
        RECT 98.710 112.155 98.880 112.615 ;
        RECT 99.550 112.155 99.720 112.615 ;
        RECT 100.390 112.155 100.560 112.615 ;
        RECT 101.230 112.155 101.535 112.615 ;
        RECT 104.620 112.155 104.895 112.975 ;
        RECT 105.565 112.155 105.735 112.625 ;
        RECT 106.405 112.155 106.575 112.625 ;
        RECT 107.245 112.155 107.415 112.625 ;
        RECT 108.085 112.155 108.255 112.625 ;
        RECT 108.925 112.155 109.095 112.625 ;
        RECT 109.765 112.155 109.935 112.625 ;
        RECT 110.605 112.155 110.775 112.625 ;
        RECT 111.445 112.155 111.735 112.625 ;
        RECT 115.535 112.155 115.865 112.635 ;
        RECT 116.375 112.155 116.705 112.635 ;
        RECT 117.215 112.155 117.545 112.635 ;
        RECT 118.055 112.155 118.385 112.635 ;
        RECT 118.895 112.155 119.225 112.635 ;
        RECT 119.735 112.155 120.065 112.955 ;
        RECT 84.530 111.985 84.990 112.155 ;
        RECT 87.030 111.985 94.390 112.155 ;
        RECT 97.530 111.985 101.670 112.155 ;
        RECT 104.530 111.985 111.890 112.155 ;
        RECT 115.020 111.985 120.540 112.155 ;
        RECT 85.605 106.665 85.895 107.390 ;
        RECT 86.915 106.665 87.085 107.145 ;
        RECT 87.755 106.665 87.925 107.145 ;
        RECT 88.595 106.665 88.765 107.145 ;
        RECT 89.435 106.665 89.605 107.145 ;
        RECT 85.520 106.495 85.980 106.665 ;
        RECT 86.320 106.495 93.680 106.665 ;
      LAYER met1 ;
        RECT 83.030 125.830 93.730 126.310 ;
        RECT 83.030 119.310 83.510 125.830 ;
        RECT 83.030 118.830 120.550 119.310 ;
        RECT 67.790 117.170 78.375 117.285 ;
        RECT 83.030 117.170 83.510 118.830 ;
        RECT 67.790 116.690 83.510 117.170 ;
        RECT 67.790 116.580 78.375 116.690 ;
        RECT 83.030 112.305 83.510 116.690 ;
        RECT 84.530 112.305 84.990 112.310 ;
        RECT 87.030 112.305 94.390 112.310 ;
        RECT 97.530 112.305 101.670 112.310 ;
        RECT 104.530 112.305 111.890 112.310 ;
        RECT 115.020 112.305 120.540 112.310 ;
        RECT 83.030 111.835 120.540 112.305 ;
        RECT 83.030 111.830 111.890 111.835 ;
        RECT 115.020 111.830 120.540 111.835 ;
        RECT 83.030 106.820 83.510 111.830 ;
        RECT 83.030 106.340 93.680 106.820 ;
      LAYER met2 ;
        RECT 46.900 117.285 59.825 117.425 ;
        RECT 67.820 117.285 68.525 117.315 ;
        RECT 46.900 116.580 68.525 117.285 ;
        RECT 46.900 116.435 59.825 116.580 ;
        RECT 67.820 116.550 68.525 116.580 ;
      LAYER met3 ;
        RECT 12.365 117.425 31.025 117.565 ;
        RECT 46.920 117.425 47.960 117.450 ;
        RECT 12.365 116.435 47.960 117.425 ;
        RECT 12.365 116.295 31.025 116.435 ;
        RECT 46.920 116.410 47.960 116.435 ;
      LAYER met4 ;
        RECT 4.000 117.565 6.000 220.760 ;
        RECT 12.390 117.565 13.670 117.570 ;
        RECT 4.000 116.295 13.670 117.565 ;
        RECT 4.000 5.000 6.000 116.295 ;
        RECT 12.390 116.290 13.670 116.295 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 86.460 126.805 90.075 126.975 ;
        RECT 86.460 126.325 86.795 126.805 ;
        RECT 87.305 126.325 87.635 126.805 ;
        RECT 88.145 126.325 88.475 126.805 ;
        RECT 88.985 126.325 89.315 126.805 ;
        RECT 89.825 126.555 90.075 126.805 ;
        RECT 93.265 126.555 93.640 126.975 ;
        RECT 89.825 126.325 93.640 126.555 ;
        RECT 98.200 120.735 98.530 121.535 ;
        RECT 99.040 120.735 99.370 121.535 ;
        RECT 99.880 120.735 100.210 121.535 ;
        RECT 100.720 120.735 101.050 121.535 ;
        RECT 104.630 120.735 104.945 121.535 ;
        RECT 105.535 120.735 105.785 121.535 ;
        RECT 106.375 120.735 106.625 121.535 ;
        RECT 107.215 120.735 107.465 121.535 ;
        RECT 108.055 121.365 111.665 121.535 ;
        RECT 108.055 120.735 108.305 121.365 ;
        RECT 97.605 120.565 101.575 120.735 ;
        RECT 91.320 120.145 93.335 120.345 ;
        RECT 97.605 119.975 97.950 120.565 ;
        RECT 101.255 119.975 101.575 120.565 ;
        RECT 104.630 120.525 108.305 120.735 ;
        RECT 108.475 120.685 108.725 121.195 ;
        RECT 108.895 120.855 109.145 121.365 ;
        RECT 109.315 120.685 109.565 121.195 ;
        RECT 109.735 120.855 109.985 121.365 ;
        RECT 110.155 120.685 110.405 121.195 ;
        RECT 110.575 120.855 110.825 121.365 ;
        RECT 110.995 120.685 111.245 121.195 ;
        RECT 111.415 120.855 111.665 121.365 ;
        RECT 115.125 120.685 115.455 121.535 ;
        RECT 115.965 120.685 116.295 121.535 ;
        RECT 108.475 120.515 111.815 120.685 ;
        RECT 115.125 120.515 116.625 120.685 ;
        RECT 104.900 120.145 108.070 120.345 ;
        RECT 108.340 120.145 111.080 120.345 ;
        RECT 111.250 119.975 111.815 120.515 ;
        RECT 115.170 120.145 116.270 120.345 ;
        RECT 116.450 120.315 116.625 120.515 ;
        RECT 116.450 120.145 119.075 120.315 ;
        RECT 116.450 119.975 116.625 120.145 ;
        RECT 87.120 119.805 90.735 119.975 ;
        RECT 87.120 119.325 87.455 119.805 ;
        RECT 87.965 119.325 88.295 119.805 ;
        RECT 88.805 119.325 89.135 119.805 ;
        RECT 89.645 119.325 89.975 119.805 ;
        RECT 90.485 119.555 90.735 119.805 ;
        RECT 93.925 119.555 94.300 119.975 ;
        RECT 97.605 119.785 101.575 119.975 ;
        RECT 105.075 119.795 111.815 119.975 ;
        RECT 115.205 119.805 116.625 119.975 ;
        RECT 90.485 119.325 94.300 119.555 ;
        RECT 98.200 119.325 98.530 119.785 ;
        RECT 99.040 119.325 99.370 119.785 ;
        RECT 99.880 119.325 100.210 119.785 ;
        RECT 100.720 119.325 101.050 119.785 ;
        RECT 105.075 119.325 105.405 119.795 ;
        RECT 105.915 119.325 106.245 119.795 ;
        RECT 106.755 119.325 107.085 119.795 ;
        RECT 107.595 119.325 107.925 119.795 ;
        RECT 108.435 119.325 108.765 119.795 ;
        RECT 109.275 119.325 109.605 119.795 ;
        RECT 110.115 119.325 110.445 119.795 ;
        RECT 110.955 119.325 111.285 119.795 ;
        RECT 115.205 119.325 115.375 119.805 ;
        RECT 116.045 119.330 116.215 119.805 ;
        RECT 98.210 113.735 98.540 114.535 ;
        RECT 99.050 113.735 99.380 114.535 ;
        RECT 99.890 113.735 100.220 114.535 ;
        RECT 100.730 113.735 101.060 114.535 ;
        RECT 104.620 113.735 104.935 114.535 ;
        RECT 105.525 113.735 105.775 114.535 ;
        RECT 106.365 113.735 106.615 114.535 ;
        RECT 107.205 113.735 107.455 114.535 ;
        RECT 108.045 114.365 111.655 114.535 ;
        RECT 108.045 113.735 108.295 114.365 ;
        RECT 97.615 113.565 101.585 113.735 ;
        RECT 87.540 113.145 90.395 113.365 ;
        RECT 97.615 112.975 97.960 113.565 ;
        RECT 101.265 112.975 101.585 113.565 ;
        RECT 104.620 113.525 108.295 113.735 ;
        RECT 108.465 113.685 108.715 114.195 ;
        RECT 108.885 113.855 109.135 114.365 ;
        RECT 109.305 113.685 109.555 114.195 ;
        RECT 109.725 113.855 109.975 114.365 ;
        RECT 110.145 113.685 110.395 114.195 ;
        RECT 110.565 113.855 110.815 114.365 ;
        RECT 110.985 113.685 111.235 114.195 ;
        RECT 111.405 113.855 111.655 114.365 ;
        RECT 115.115 113.685 115.445 114.535 ;
        RECT 115.955 113.685 116.285 114.535 ;
        RECT 108.465 113.515 111.805 113.685 ;
        RECT 115.115 113.515 116.615 113.685 ;
        RECT 104.890 113.145 108.060 113.345 ;
        RECT 108.330 113.145 111.070 113.345 ;
        RECT 111.240 112.975 111.805 113.515 ;
        RECT 115.160 113.145 116.260 113.345 ;
        RECT 116.440 113.315 116.615 113.515 ;
        RECT 116.440 113.145 119.065 113.315 ;
        RECT 116.440 112.975 116.615 113.145 ;
        RECT 87.120 112.805 90.735 112.975 ;
        RECT 87.120 112.325 87.455 112.805 ;
        RECT 87.965 112.325 88.295 112.805 ;
        RECT 88.805 112.325 89.135 112.805 ;
        RECT 89.645 112.325 89.975 112.805 ;
        RECT 90.485 112.555 90.735 112.805 ;
        RECT 93.925 112.555 94.300 112.975 ;
        RECT 97.615 112.785 101.585 112.975 ;
        RECT 105.065 112.795 111.805 112.975 ;
        RECT 115.195 112.805 116.615 112.975 ;
        RECT 90.485 112.325 94.300 112.555 ;
        RECT 98.210 112.325 98.540 112.785 ;
        RECT 99.050 112.325 99.380 112.785 ;
        RECT 99.890 112.325 100.220 112.785 ;
        RECT 100.730 112.325 101.060 112.785 ;
        RECT 105.065 112.325 105.395 112.795 ;
        RECT 105.905 112.325 106.235 112.795 ;
        RECT 106.745 112.325 107.075 112.795 ;
        RECT 107.585 112.325 107.915 112.795 ;
        RECT 108.425 112.325 108.755 112.795 ;
        RECT 109.265 112.325 109.595 112.795 ;
        RECT 110.105 112.325 110.435 112.795 ;
        RECT 110.945 112.325 111.275 112.795 ;
        RECT 115.195 112.325 115.365 112.805 ;
        RECT 116.035 112.330 116.205 112.805 ;
        RECT 86.410 107.315 90.025 107.485 ;
        RECT 86.410 106.835 86.745 107.315 ;
        RECT 87.255 106.835 87.585 107.315 ;
        RECT 88.095 106.835 88.425 107.315 ;
        RECT 88.935 106.835 89.265 107.315 ;
        RECT 89.775 107.065 90.025 107.315 ;
        RECT 93.215 107.065 93.590 107.485 ;
        RECT 89.775 106.835 93.590 107.065 ;
      LAYER met1 ;
        RECT 92.740 120.030 93.190 120.450 ;
        RECT 101.270 120.350 101.560 120.365 ;
        RECT 105.450 120.350 105.870 120.410 ;
        RECT 101.270 120.145 105.870 120.350 ;
        RECT 101.270 120.135 101.560 120.145 ;
        RECT 105.450 120.080 105.870 120.145 ;
        RECT 108.850 120.030 109.190 120.410 ;
        RECT 111.460 120.310 111.750 120.340 ;
        RECT 112.565 120.310 112.885 120.350 ;
        RECT 115.330 120.310 115.670 120.430 ;
        RECT 111.460 120.135 115.670 120.310 ;
        RECT 111.460 120.110 111.750 120.135 ;
        RECT 112.565 120.090 112.885 120.135 ;
        RECT 115.330 120.030 115.670 120.135 ;
        RECT 92.845 119.820 93.075 120.030 ;
        RECT 108.940 119.830 109.110 120.030 ;
        RECT 92.830 119.500 93.090 119.820 ;
        RECT 108.895 119.510 109.155 119.830 ;
        RECT 92.800 118.115 93.120 118.130 ;
        RECT 110.260 118.115 110.580 118.130 ;
        RECT 92.800 117.885 110.580 118.115 ;
        RECT 92.800 117.870 93.120 117.885 ;
        RECT 110.260 117.870 110.580 117.885 ;
        RECT 113.275 115.965 113.595 115.990 ;
        RECT 89.040 115.760 113.595 115.965 ;
        RECT 89.040 115.570 89.245 115.760 ;
        RECT 113.275 115.730 113.595 115.760 ;
        RECT 88.980 115.310 89.300 115.570 ;
        RECT 89.005 113.840 89.265 114.160 ;
        RECT 111.360 113.970 111.680 114.230 ;
        RECT 89.030 113.430 89.235 113.840 ;
        RECT 103.425 113.740 108.760 113.910 ;
        RECT 88.960 113.100 89.270 113.430 ;
        RECT 101.305 113.315 101.595 113.345 ;
        RECT 103.425 113.315 103.595 113.740 ;
        RECT 108.590 113.420 108.760 113.740 ;
        RECT 101.305 113.145 103.595 113.315 ;
        RECT 101.305 113.115 101.595 113.145 ;
        RECT 106.120 113.030 106.500 113.410 ;
        RECT 108.520 113.090 108.820 113.420 ;
        RECT 111.435 113.365 111.605 113.970 ;
        RECT 113.300 113.800 113.560 114.120 ;
        RECT 111.405 113.350 111.635 113.365 ;
        RECT 113.325 113.350 113.530 113.800 ;
        RECT 115.340 113.350 115.670 113.420 ;
        RECT 111.405 113.145 115.670 113.350 ;
        RECT 111.405 113.075 111.635 113.145 ;
        RECT 115.340 113.080 115.670 113.145 ;
        RECT 106.235 112.750 106.410 113.030 ;
        RECT 112.560 112.750 112.880 112.795 ;
        RECT 106.235 112.575 112.880 112.750 ;
        RECT 106.235 112.560 106.410 112.575 ;
        RECT 112.560 112.535 112.880 112.575 ;
      LAYER met2 ;
        RECT 112.595 120.060 112.855 120.380 ;
        RECT 92.800 119.530 93.120 119.790 ;
        RECT 108.865 119.540 109.185 119.800 ;
        RECT 92.845 118.160 93.075 119.530 ;
        RECT 92.830 117.840 93.090 118.160 ;
        RECT 108.940 116.365 109.110 119.540 ;
        RECT 110.290 118.115 110.550 118.160 ;
        RECT 112.635 118.115 112.810 120.060 ;
        RECT 110.290 117.885 112.810 118.115 ;
        RECT 110.290 117.840 110.550 117.885 ;
        RECT 108.940 116.195 111.605 116.365 ;
        RECT 89.010 115.280 89.270 115.600 ;
        RECT 89.035 114.130 89.240 115.280 ;
        RECT 111.435 114.260 111.605 116.195 ;
        RECT 88.975 113.870 89.295 114.130 ;
        RECT 111.390 113.940 111.650 114.260 ;
        RECT 112.635 112.825 112.810 117.885 ;
        RECT 113.305 115.700 113.565 116.020 ;
        RECT 113.330 114.090 113.535 115.700 ;
        RECT 113.270 113.830 113.590 114.090 ;
        RECT 112.590 112.505 112.850 112.825 ;
  END
END tt_um_relax
END LIBRARY

