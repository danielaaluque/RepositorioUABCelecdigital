VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO layout
  CLASS BLOCK ;
  FOREIGN layout ;
  ORIGIN 19.680 16.380 ;
  SIZE 44.850 BY 26.500 ;
  OBS
      LAYER pwell ;
        RECT -9.730 9.485 -8.945 9.915 ;
      LAYER nwell ;
        RECT -8.615 9.280 -7.010 10.120 ;
        RECT -8.150 6.780 -7.310 9.280 ;
        RECT -12.680 5.175 -4.940 6.780 ;
      LAYER pwell ;
        RECT -12.485 3.975 -5.135 4.885 ;
        RECT -12.340 3.785 -12.170 3.975 ;
        RECT -1.410 3.225 -0.625 3.655 ;
      LAYER nwell ;
        RECT -0.295 3.020 1.310 3.860 ;
      LAYER pwell ;
        RECT 7.020 3.225 7.805 3.655 ;
      LAYER nwell ;
        RECT 8.135 3.020 9.740 3.860 ;
        RECT 0.060 0.950 0.900 3.020 ;
        RECT -14.170 -0.715 -4.780 0.890 ;
        RECT -3.350 -0.655 1.170 0.950 ;
        RECT 8.520 0.670 9.360 3.020 ;
      LAYER pwell ;
        RECT -13.975 -1.915 -6.625 -1.005 ;
        RECT -13.830 -2.105 -13.660 -1.915 ;
      LAYER nwell ;
        RECT -6.385 -2.655 -4.780 -0.715 ;
        RECT 4.430 -0.935 12.170 0.670 ;
      LAYER pwell ;
        RECT -2.990 -1.855 0.880 -0.945 ;
      LAYER nwell ;
        RECT 14.640 -1.005 22.760 0.600 ;
      LAYER pwell ;
        RECT -2.990 -1.875 -2.845 -1.855 ;
        RECT -3.015 -2.045 -2.845 -1.875 ;
        RECT 4.625 -2.135 11.875 -1.225 ;
        RECT 4.765 -2.325 4.935 -2.135 ;
        RECT 14.835 -2.205 19.965 -1.295 ;
        RECT 22.125 -2.120 22.555 -1.335 ;
        RECT 14.980 -2.395 15.150 -2.205 ;
      LAYER nwell ;
        RECT -9.480 -3.210 -4.780 -2.655 ;
      LAYER pwell ;
        RECT -11.600 -3.845 -10.815 -3.415 ;
      LAYER nwell ;
        RECT -10.485 -4.050 -4.780 -3.210 ;
        RECT -9.480 -4.260 -4.780 -4.050 ;
      LAYER pwell ;
        RECT 5.570 -5.335 6.355 -4.905 ;
      LAYER nwell ;
        RECT 6.685 -5.540 8.290 -4.700 ;
        RECT -19.680 -7.210 -18.840 -7.040 ;
        RECT -19.680 -8.645 -6.150 -7.210 ;
        RECT 7.050 -7.220 7.890 -5.540 ;
        RECT -19.060 -8.815 -6.150 -8.645 ;
        RECT -3.460 -8.825 2.610 -7.220 ;
        RECT 4.430 -8.825 12.170 -7.220 ;
        RECT 14.390 -7.390 22.610 -7.350 ;
      LAYER pwell ;
        RECT -19.475 -9.760 -19.045 -8.975 ;
        RECT -13.695 -10.015 -6.345 -9.105 ;
        RECT -13.550 -10.205 -13.380 -10.015 ;
        RECT -3.100 -10.025 0.770 -9.115 ;
        RECT -3.100 -10.045 -2.955 -10.025 ;
        RECT -3.125 -10.215 -2.955 -10.045 ;
      LAYER nwell ;
        RECT 1.005 -11.060 2.610 -8.825 ;
        RECT 14.390 -8.955 23.240 -7.390 ;
        RECT 22.400 -8.995 23.240 -8.955 ;
      LAYER pwell ;
        RECT 4.625 -10.025 11.875 -9.115 ;
        RECT 4.765 -10.215 4.935 -10.025 ;
        RECT 14.585 -10.155 19.715 -9.245 ;
        RECT 22.605 -10.110 23.035 -9.325 ;
        RECT 14.730 -10.345 14.900 -10.155 ;
        RECT -1.400 -11.695 -0.615 -11.265 ;
      LAYER nwell ;
        RECT -0.285 -11.900 2.610 -11.060 ;
        RECT 1.005 -11.930 2.610 -11.900 ;
        RECT -2.420 -12.870 -1.580 -12.640 ;
        RECT -13.000 -14.245 -1.580 -12.870 ;
        RECT -13.000 -14.475 -2.020 -14.245 ;
      LAYER pwell ;
        RECT -12.805 -15.675 -5.455 -14.765 ;
        RECT -2.215 -15.360 -1.785 -14.575 ;
        RECT -12.660 -15.865 -12.490 -15.675 ;
      LAYER li1 ;
        RECT -10.005 9.845 -9.835 9.930 ;
        RECT -7.285 9.845 -7.115 9.930 ;
        RECT -10.005 9.555 -9.110 9.845 ;
        RECT -8.450 9.555 -7.115 9.845 ;
        RECT -10.005 9.470 -9.835 9.555 ;
        RECT -7.285 9.470 -7.115 9.555 ;
        RECT -12.490 6.505 -5.130 6.675 ;
        RECT -12.400 5.365 -12.145 6.505 ;
        RECT -11.975 5.535 -11.645 6.335 ;
        RECT -11.475 5.705 -11.305 6.505 ;
        RECT -11.135 5.535 -10.805 6.335 ;
        RECT -10.635 5.705 -10.465 6.505 ;
        RECT -10.295 5.535 -9.965 6.335 ;
        RECT -9.795 5.705 -9.625 6.505 ;
        RECT -9.455 5.535 -9.125 6.335 ;
        RECT -8.955 5.705 -8.785 6.505 ;
        RECT -8.615 5.535 -8.285 6.335 ;
        RECT -8.115 5.705 -7.945 6.505 ;
        RECT -7.775 5.535 -7.445 6.335 ;
        RECT -7.275 5.705 -7.105 6.505 ;
        RECT -6.935 5.535 -6.605 6.335 ;
        RECT -6.435 5.705 -6.265 6.505 ;
        RECT -6.095 5.535 -5.765 6.335 ;
        RECT -11.975 5.335 -5.765 5.535 ;
        RECT -5.575 5.365 -5.220 6.505 ;
        RECT -11.980 4.945 -9.125 5.165 ;
        RECT -8.850 4.945 -8.370 5.335 ;
        RECT -8.200 4.945 -6.185 5.145 ;
        RECT -8.615 4.775 -8.370 4.945 ;
        RECT -6.015 4.775 -5.765 5.335 ;
        RECT -12.400 4.605 -8.785 4.775 ;
        RECT -12.400 4.125 -12.065 4.605 ;
        RECT -11.895 3.955 -11.725 4.435 ;
        RECT -11.555 4.125 -11.225 4.605 ;
        RECT -11.055 3.955 -10.885 4.435 ;
        RECT -10.715 4.125 -10.385 4.605 ;
        RECT -10.215 3.955 -10.045 4.435 ;
        RECT -9.875 4.125 -9.545 4.605 ;
        RECT -9.375 3.955 -9.205 4.435 ;
        RECT -9.035 4.355 -8.785 4.605 ;
        RECT -8.615 4.525 -5.765 4.775 ;
        RECT -5.595 4.355 -5.220 4.775 ;
        RECT -9.035 4.125 -5.220 4.355 ;
        RECT -12.490 3.785 -5.130 3.955 ;
        RECT -1.685 3.585 -1.515 3.670 ;
        RECT 1.035 3.585 1.205 3.670 ;
        RECT -1.685 3.295 -0.790 3.585 ;
        RECT -0.130 3.295 1.205 3.585 ;
        RECT -1.685 3.210 -1.515 3.295 ;
        RECT 1.035 3.210 1.205 3.295 ;
        RECT 6.745 3.585 6.915 3.670 ;
        RECT 9.465 3.585 9.635 3.670 ;
        RECT 6.745 3.295 7.640 3.585 ;
        RECT 8.300 3.295 9.635 3.585 ;
        RECT 6.745 3.210 6.915 3.295 ;
        RECT 9.465 3.210 9.635 3.295 ;
        RECT -13.980 0.615 -6.620 0.785 ;
        RECT -3.160 0.675 0.980 0.845 ;
        RECT -13.890 -0.525 -13.635 0.615 ;
        RECT -13.465 -0.355 -13.135 0.445 ;
        RECT -12.965 -0.185 -12.795 0.615 ;
        RECT -12.625 -0.355 -12.295 0.445 ;
        RECT -12.125 -0.185 -11.955 0.615 ;
        RECT -11.785 -0.355 -11.455 0.445 ;
        RECT -11.285 -0.185 -11.115 0.615 ;
        RECT -10.945 -0.355 -10.615 0.445 ;
        RECT -10.445 -0.185 -10.275 0.615 ;
        RECT -10.105 -0.355 -9.775 0.445 ;
        RECT -9.605 -0.185 -9.435 0.615 ;
        RECT -9.265 -0.355 -8.935 0.445 ;
        RECT -8.765 -0.185 -8.595 0.615 ;
        RECT -8.425 -0.355 -8.095 0.445 ;
        RECT -7.925 -0.185 -7.755 0.615 ;
        RECT -7.585 -0.355 -7.255 0.445 ;
        RECT -13.465 -0.555 -7.255 -0.355 ;
        RECT -7.065 -0.525 -6.710 0.615 ;
        RECT -2.905 -0.125 -2.650 0.675 ;
        RECT -2.480 -0.295 -2.150 0.505 ;
        RECT -1.980 -0.125 -1.810 0.675 ;
        RECT -1.640 -0.295 -1.310 0.505 ;
        RECT -1.140 -0.125 -0.970 0.675 ;
        RECT -0.800 -0.295 -0.470 0.505 ;
        RECT -0.300 -0.125 -0.130 0.675 ;
        RECT 0.040 -0.295 0.370 0.505 ;
        RECT 0.540 -0.125 0.840 0.675 ;
        RECT 4.620 0.395 11.980 0.565 ;
        RECT -3.075 -0.465 0.895 -0.295 ;
        RECT -13.470 -0.945 -10.615 -0.725 ;
        RECT -10.340 -0.945 -9.860 -0.555 ;
        RECT -9.690 -0.945 -7.675 -0.745 ;
        RECT -10.105 -1.115 -9.860 -0.945 ;
        RECT -7.505 -1.115 -7.255 -0.555 ;
        RECT -3.075 -1.055 -2.730 -0.465 ;
        RECT -2.480 -0.885 0.375 -0.635 ;
        RECT 0.575 -1.055 0.895 -0.465 ;
        RECT 4.710 -0.575 5.025 0.225 ;
        RECT 5.195 -0.405 5.445 0.395 ;
        RECT 5.615 -0.575 5.865 0.225 ;
        RECT 6.035 -0.405 6.285 0.395 ;
        RECT 6.455 -0.575 6.705 0.225 ;
        RECT 6.875 -0.405 7.125 0.395 ;
        RECT 7.295 -0.575 7.545 0.225 ;
        RECT 7.715 -0.405 7.965 0.395 ;
        RECT 14.830 0.325 20.350 0.495 ;
        RECT 22.110 0.325 22.570 0.495 ;
        RECT 8.135 0.055 11.745 0.225 ;
        RECT 8.135 -0.575 8.385 0.055 ;
        RECT 4.710 -0.785 8.385 -0.575 ;
        RECT 8.555 -0.625 8.805 -0.115 ;
        RECT 8.975 -0.455 9.225 0.055 ;
        RECT 9.395 -0.625 9.645 -0.115 ;
        RECT 9.815 -0.455 10.065 0.055 ;
        RECT 10.235 -0.625 10.485 -0.115 ;
        RECT 10.655 -0.455 10.905 0.055 ;
        RECT 11.075 -0.625 11.325 -0.115 ;
        RECT 11.495 -0.455 11.745 0.055 ;
        RECT 8.555 -0.795 11.895 -0.625 ;
        RECT -13.890 -1.285 -10.275 -1.115 ;
        RECT -13.890 -1.765 -13.555 -1.285 ;
        RECT -13.385 -1.935 -13.215 -1.455 ;
        RECT -13.045 -1.765 -12.715 -1.285 ;
        RECT -12.545 -1.935 -12.375 -1.455 ;
        RECT -12.205 -1.765 -11.875 -1.285 ;
        RECT -11.705 -1.935 -11.535 -1.455 ;
        RECT -11.365 -1.765 -11.035 -1.285 ;
        RECT -10.865 -1.935 -10.695 -1.455 ;
        RECT -10.525 -1.535 -10.275 -1.285 ;
        RECT -10.105 -1.365 -7.255 -1.115 ;
        RECT -7.085 -1.535 -6.710 -1.115 ;
        RECT -3.075 -1.245 0.895 -1.055 ;
        RECT 4.980 -1.165 8.150 -0.965 ;
        RECT 8.420 -1.165 11.160 -0.965 ;
        RECT -10.525 -1.765 -6.710 -1.535 ;
        RECT -2.905 -1.875 -2.650 -1.415 ;
        RECT -2.480 -1.705 -2.150 -1.245 ;
        RECT -1.980 -1.875 -1.810 -1.415 ;
        RECT -1.640 -1.705 -1.310 -1.245 ;
        RECT -1.140 -1.875 -0.970 -1.415 ;
        RECT -0.800 -1.705 -0.470 -1.245 ;
        RECT -0.300 -1.875 -0.130 -1.415 ;
        RECT 0.040 -1.705 0.370 -1.245 ;
        RECT 11.330 -1.335 11.895 -0.795 ;
        RECT 14.925 -0.695 15.255 0.155 ;
        RECT 15.425 -0.475 15.595 0.325 ;
        RECT 15.765 -0.695 16.095 0.155 ;
        RECT 16.265 -0.475 16.435 0.325 ;
        RECT 16.685 -0.695 16.855 0.155 ;
        RECT 17.025 -0.475 17.355 0.325 ;
        RECT 17.525 -0.695 17.695 0.155 ;
        RECT 17.865 -0.475 18.195 0.325 ;
        RECT 18.365 -0.695 18.535 0.155 ;
        RECT 18.705 -0.475 19.035 0.325 ;
        RECT 19.205 -0.695 19.375 0.155 ;
        RECT 14.925 -0.865 16.425 -0.695 ;
        RECT 16.685 -0.865 19.375 -0.695 ;
        RECT 19.545 -0.825 19.875 0.325 ;
        RECT 22.195 -0.840 22.485 0.325 ;
        RECT 14.970 -1.235 16.070 -1.035 ;
        RECT 16.250 -1.065 16.425 -0.865 ;
        RECT 16.250 -1.235 18.875 -1.065 ;
        RECT 0.540 -1.875 0.845 -1.415 ;
        RECT -13.980 -2.105 -6.620 -1.935 ;
        RECT -3.160 -2.045 0.980 -1.875 ;
        RECT 4.710 -2.155 4.985 -1.335 ;
        RECT 5.155 -1.515 11.895 -1.335 ;
        RECT 16.250 -1.405 16.425 -1.235 ;
        RECT 19.120 -1.405 19.375 -0.865 ;
        RECT 5.155 -1.985 5.485 -1.515 ;
        RECT 5.655 -2.155 5.825 -1.685 ;
        RECT 5.995 -1.985 6.325 -1.515 ;
        RECT 6.495 -2.155 6.665 -1.685 ;
        RECT 6.835 -1.985 7.165 -1.515 ;
        RECT 7.335 -2.155 7.505 -1.685 ;
        RECT 7.675 -1.985 8.005 -1.515 ;
        RECT 8.175 -2.155 8.345 -1.685 ;
        RECT 8.515 -1.985 8.845 -1.515 ;
        RECT 9.015 -2.155 9.185 -1.685 ;
        RECT 9.355 -1.985 9.685 -1.515 ;
        RECT 9.855 -2.155 10.025 -1.685 ;
        RECT 10.195 -1.985 10.525 -1.515 ;
        RECT 10.695 -2.155 10.865 -1.685 ;
        RECT 11.035 -1.985 11.365 -1.515 ;
        RECT 15.005 -1.575 16.425 -1.405 ;
        RECT 16.685 -1.575 19.375 -1.405 ;
        RECT 11.535 -2.155 11.825 -1.685 ;
        RECT 15.005 -2.055 15.175 -1.575 ;
        RECT 4.620 -2.325 11.980 -2.155 ;
        RECT 15.345 -2.225 15.675 -1.745 ;
        RECT 15.845 -2.050 16.015 -1.575 ;
        RECT 16.185 -2.225 16.515 -1.745 ;
        RECT 16.685 -2.055 16.855 -1.575 ;
        RECT 17.025 -2.225 17.355 -1.745 ;
        RECT 17.525 -2.055 17.695 -1.575 ;
        RECT 17.865 -2.225 18.195 -1.745 ;
        RECT 18.365 -2.055 18.535 -1.575 ;
        RECT 18.705 -2.225 19.035 -1.745 ;
        RECT 19.205 -2.055 19.375 -1.575 ;
        RECT 19.545 -2.225 19.875 -1.425 ;
        RECT 22.195 -2.225 22.485 -1.500 ;
        RECT 14.830 -2.395 20.350 -2.225 ;
        RECT 22.110 -2.395 22.570 -2.225 ;
        RECT -11.875 -3.485 -11.705 -3.400 ;
        RECT -9.155 -3.485 -8.985 -3.400 ;
        RECT -11.875 -3.775 -10.980 -3.485 ;
        RECT -10.320 -3.775 -8.985 -3.485 ;
        RECT -11.875 -3.860 -11.705 -3.775 ;
        RECT -9.155 -3.860 -8.985 -3.775 ;
        RECT 5.295 -4.975 5.465 -4.890 ;
        RECT 8.015 -4.975 8.185 -4.890 ;
        RECT 5.295 -5.265 6.190 -4.975 ;
        RECT 6.850 -5.265 8.185 -4.975 ;
        RECT 5.295 -5.350 5.465 -5.265 ;
        RECT 8.015 -5.350 8.185 -5.265 ;
        RECT -19.490 -7.315 -19.030 -7.145 ;
        RECT -19.405 -8.480 -19.115 -7.315 ;
        RECT -13.700 -7.485 -6.340 -7.315 ;
        RECT -13.610 -8.625 -13.355 -7.485 ;
        RECT -13.185 -8.455 -12.855 -7.655 ;
        RECT -12.685 -8.285 -12.515 -7.485 ;
        RECT -12.345 -8.455 -12.015 -7.655 ;
        RECT -11.845 -8.285 -11.675 -7.485 ;
        RECT -11.505 -8.455 -11.175 -7.655 ;
        RECT -11.005 -8.285 -10.835 -7.485 ;
        RECT -10.665 -8.455 -10.335 -7.655 ;
        RECT -10.165 -8.285 -9.995 -7.485 ;
        RECT -9.825 -8.455 -9.495 -7.655 ;
        RECT -9.325 -8.285 -9.155 -7.485 ;
        RECT -8.985 -8.455 -8.655 -7.655 ;
        RECT -8.485 -8.285 -8.315 -7.485 ;
        RECT -8.145 -8.455 -7.815 -7.655 ;
        RECT -7.645 -8.285 -7.475 -7.485 ;
        RECT -7.305 -8.455 -6.975 -7.655 ;
        RECT -13.185 -8.655 -6.975 -8.455 ;
        RECT -6.785 -8.625 -6.430 -7.485 ;
        RECT -3.270 -7.495 0.870 -7.325 ;
        RECT 4.620 -7.495 11.980 -7.325 ;
        RECT -3.015 -8.295 -2.760 -7.495 ;
        RECT -2.590 -8.465 -2.260 -7.665 ;
        RECT -2.090 -8.295 -1.920 -7.495 ;
        RECT -1.750 -8.465 -1.420 -7.665 ;
        RECT -1.250 -8.295 -1.080 -7.495 ;
        RECT -0.910 -8.465 -0.580 -7.665 ;
        RECT -0.410 -8.295 -0.240 -7.495 ;
        RECT -0.070 -8.465 0.260 -7.665 ;
        RECT 0.430 -8.295 0.730 -7.495 ;
        RECT 4.710 -8.465 5.025 -7.665 ;
        RECT 5.195 -8.295 5.445 -7.495 ;
        RECT 5.615 -8.465 5.865 -7.665 ;
        RECT 6.035 -8.295 6.285 -7.495 ;
        RECT 6.455 -8.465 6.705 -7.665 ;
        RECT 6.875 -8.295 7.125 -7.495 ;
        RECT 7.295 -8.465 7.545 -7.665 ;
        RECT 7.715 -8.295 7.965 -7.495 ;
        RECT 14.580 -7.625 20.100 -7.455 ;
        RECT 8.135 -7.835 11.745 -7.665 ;
        RECT 8.135 -8.465 8.385 -7.835 ;
        RECT -13.190 -9.045 -10.335 -8.825 ;
        RECT -10.060 -9.045 -9.580 -8.655 ;
        RECT -9.410 -9.045 -7.395 -8.845 ;
        RECT -19.405 -9.865 -19.115 -9.140 ;
        RECT -9.825 -9.215 -9.580 -9.045 ;
        RECT -7.225 -9.215 -6.975 -8.655 ;
        RECT -3.185 -8.635 0.785 -8.465 ;
        RECT -13.610 -9.385 -9.995 -9.215 ;
        RECT -13.610 -9.865 -13.275 -9.385 ;
        RECT -19.490 -10.035 -19.030 -9.865 ;
        RECT -13.105 -10.035 -12.935 -9.555 ;
        RECT -12.765 -9.865 -12.435 -9.385 ;
        RECT -12.265 -10.035 -12.095 -9.555 ;
        RECT -11.925 -9.865 -11.595 -9.385 ;
        RECT -11.425 -10.035 -11.255 -9.555 ;
        RECT -11.085 -9.865 -10.755 -9.385 ;
        RECT -10.585 -10.035 -10.415 -9.555 ;
        RECT -10.245 -9.635 -9.995 -9.385 ;
        RECT -9.825 -9.465 -6.975 -9.215 ;
        RECT -6.805 -9.635 -6.430 -9.215 ;
        RECT -3.185 -9.225 -2.840 -8.635 ;
        RECT -2.590 -9.055 0.265 -8.805 ;
        RECT 0.465 -9.225 0.785 -8.635 ;
        RECT 4.710 -8.675 8.385 -8.465 ;
        RECT 8.555 -8.515 8.805 -8.005 ;
        RECT 8.975 -8.345 9.225 -7.835 ;
        RECT 9.395 -8.515 9.645 -8.005 ;
        RECT 9.815 -8.345 10.065 -7.835 ;
        RECT 10.235 -8.515 10.485 -8.005 ;
        RECT 10.655 -8.345 10.905 -7.835 ;
        RECT 11.075 -8.515 11.325 -8.005 ;
        RECT 11.495 -8.345 11.745 -7.835 ;
        RECT 8.555 -8.685 11.895 -8.515 ;
        RECT 4.980 -9.055 8.150 -8.855 ;
        RECT 8.420 -9.055 11.160 -8.855 ;
        RECT 11.330 -9.225 11.895 -8.685 ;
        RECT 14.675 -8.645 15.005 -7.795 ;
        RECT 15.175 -8.425 15.345 -7.625 ;
        RECT 15.515 -8.645 15.845 -7.795 ;
        RECT 16.015 -8.425 16.185 -7.625 ;
        RECT 16.435 -8.645 16.605 -7.795 ;
        RECT 16.775 -8.425 17.105 -7.625 ;
        RECT 17.275 -8.645 17.445 -7.795 ;
        RECT 17.615 -8.425 17.945 -7.625 ;
        RECT 18.115 -8.645 18.285 -7.795 ;
        RECT 18.455 -8.425 18.785 -7.625 ;
        RECT 18.955 -8.645 19.125 -7.795 ;
        RECT 14.675 -8.815 16.175 -8.645 ;
        RECT 16.435 -8.815 19.125 -8.645 ;
        RECT 19.295 -8.775 19.625 -7.625 ;
        RECT 22.590 -7.665 23.050 -7.495 ;
        RECT 14.720 -9.185 15.820 -8.985 ;
        RECT 16.000 -9.015 16.175 -8.815 ;
        RECT 16.000 -9.185 18.625 -9.015 ;
        RECT -3.185 -9.415 0.785 -9.225 ;
        RECT -10.245 -9.865 -6.430 -9.635 ;
        RECT -13.700 -10.205 -6.340 -10.035 ;
        RECT -3.015 -10.045 -2.760 -9.585 ;
        RECT -2.590 -9.875 -2.260 -9.415 ;
        RECT -2.090 -10.045 -1.920 -9.585 ;
        RECT -1.750 -9.875 -1.420 -9.415 ;
        RECT -1.250 -10.045 -1.080 -9.585 ;
        RECT -0.910 -9.875 -0.580 -9.415 ;
        RECT -0.410 -10.045 -0.240 -9.585 ;
        RECT -0.070 -9.875 0.260 -9.415 ;
        RECT 0.430 -10.045 0.735 -9.585 ;
        RECT 4.710 -10.045 4.985 -9.225 ;
        RECT 5.155 -9.405 11.895 -9.225 ;
        RECT 16.000 -9.355 16.175 -9.185 ;
        RECT 18.870 -9.355 19.125 -8.815 ;
        RECT 22.675 -8.830 22.965 -7.665 ;
        RECT 5.155 -9.875 5.485 -9.405 ;
        RECT 5.655 -10.045 5.825 -9.575 ;
        RECT 5.995 -9.875 6.325 -9.405 ;
        RECT 6.495 -10.045 6.665 -9.575 ;
        RECT 6.835 -9.875 7.165 -9.405 ;
        RECT 7.335 -10.045 7.505 -9.575 ;
        RECT 7.675 -9.875 8.005 -9.405 ;
        RECT 8.175 -10.045 8.345 -9.575 ;
        RECT 8.515 -9.875 8.845 -9.405 ;
        RECT 9.015 -10.045 9.185 -9.575 ;
        RECT 9.355 -9.875 9.685 -9.405 ;
        RECT 9.855 -10.045 10.025 -9.575 ;
        RECT 10.195 -9.875 10.525 -9.405 ;
        RECT 10.695 -10.045 10.865 -9.575 ;
        RECT 11.035 -9.875 11.365 -9.405 ;
        RECT 14.755 -9.525 16.175 -9.355 ;
        RECT 16.435 -9.525 19.125 -9.355 ;
        RECT 11.535 -10.045 11.825 -9.575 ;
        RECT 14.755 -10.005 14.925 -9.525 ;
        RECT -3.270 -10.215 0.870 -10.045 ;
        RECT 4.620 -10.215 11.980 -10.045 ;
        RECT 15.095 -10.175 15.425 -9.695 ;
        RECT 15.595 -10.000 15.765 -9.525 ;
        RECT 15.935 -10.175 16.265 -9.695 ;
        RECT 16.435 -10.005 16.605 -9.525 ;
        RECT 16.775 -10.175 17.105 -9.695 ;
        RECT 17.275 -10.005 17.445 -9.525 ;
        RECT 17.615 -10.175 17.945 -9.695 ;
        RECT 18.115 -10.005 18.285 -9.525 ;
        RECT 18.455 -10.175 18.785 -9.695 ;
        RECT 18.955 -10.005 19.125 -9.525 ;
        RECT 19.295 -10.175 19.625 -9.375 ;
        RECT 14.580 -10.345 20.100 -10.175 ;
        RECT 22.675 -10.215 22.965 -9.490 ;
        RECT 22.590 -10.385 23.050 -10.215 ;
        RECT -1.675 -11.335 -1.505 -11.250 ;
        RECT 1.045 -11.335 1.215 -11.250 ;
        RECT -1.675 -11.625 -0.780 -11.335 ;
        RECT -0.120 -11.625 1.215 -11.335 ;
        RECT -1.675 -11.710 -1.505 -11.625 ;
        RECT 1.045 -11.710 1.215 -11.625 ;
        RECT -2.230 -12.915 -1.770 -12.745 ;
        RECT -12.810 -13.145 -5.450 -12.975 ;
        RECT -12.720 -14.285 -12.465 -13.145 ;
        RECT -12.295 -14.115 -11.965 -13.315 ;
        RECT -11.795 -13.945 -11.625 -13.145 ;
        RECT -11.455 -14.115 -11.125 -13.315 ;
        RECT -10.955 -13.945 -10.785 -13.145 ;
        RECT -10.615 -14.115 -10.285 -13.315 ;
        RECT -10.115 -13.945 -9.945 -13.145 ;
        RECT -9.775 -14.115 -9.445 -13.315 ;
        RECT -9.275 -13.945 -9.105 -13.145 ;
        RECT -8.935 -14.115 -8.605 -13.315 ;
        RECT -8.435 -13.945 -8.265 -13.145 ;
        RECT -8.095 -14.115 -7.765 -13.315 ;
        RECT -7.595 -13.945 -7.425 -13.145 ;
        RECT -7.255 -14.115 -6.925 -13.315 ;
        RECT -6.755 -13.945 -6.585 -13.145 ;
        RECT -6.415 -14.115 -6.085 -13.315 ;
        RECT -12.295 -14.315 -6.085 -14.115 ;
        RECT -5.895 -14.285 -5.540 -13.145 ;
        RECT -2.145 -14.080 -1.855 -12.915 ;
        RECT -12.300 -14.705 -9.445 -14.485 ;
        RECT -9.170 -14.705 -8.690 -14.315 ;
        RECT -8.520 -14.705 -6.505 -14.505 ;
        RECT -8.935 -14.875 -8.690 -14.705 ;
        RECT -6.335 -14.875 -6.085 -14.315 ;
        RECT -12.720 -15.045 -9.105 -14.875 ;
        RECT -12.720 -15.525 -12.385 -15.045 ;
        RECT -12.215 -15.695 -12.045 -15.215 ;
        RECT -11.875 -15.525 -11.545 -15.045 ;
        RECT -11.375 -15.695 -11.205 -15.215 ;
        RECT -11.035 -15.525 -10.705 -15.045 ;
        RECT -10.535 -15.695 -10.365 -15.215 ;
        RECT -10.195 -15.525 -9.865 -15.045 ;
        RECT -9.695 -15.695 -9.525 -15.215 ;
        RECT -9.355 -15.295 -9.105 -15.045 ;
        RECT -8.935 -15.125 -6.085 -14.875 ;
        RECT -5.915 -15.295 -5.540 -14.875 ;
        RECT -9.355 -15.525 -5.540 -15.295 ;
        RECT -2.145 -15.465 -1.855 -14.740 ;
        RECT -2.230 -15.635 -1.770 -15.465 ;
        RECT -12.810 -15.865 -5.450 -15.695 ;
      LAYER met1 ;
        RECT -10.160 9.470 -9.680 9.930 ;
        RECT -7.440 9.470 -6.960 9.930 ;
        RECT -10.160 7.955 -10.005 9.470 ;
        RECT -10.240 7.695 -9.920 7.955 ;
        RECT -14.725 6.830 -14.435 6.860 ;
        RECT -7.115 6.830 -6.960 9.470 ;
        RECT -14.725 6.675 2.125 6.830 ;
        RECT -14.725 6.540 -5.130 6.675 ;
        RECT -14.725 6.510 -14.435 6.540 ;
        RECT -12.490 6.350 -5.130 6.540 ;
        RECT -9.020 5.430 -8.170 5.530 ;
        RECT -11.730 5.165 -11.450 5.195 ;
        RECT -13.180 4.945 -11.060 5.165 ;
        RECT -9.020 5.050 -2.830 5.430 ;
        RECT -1.180 5.290 -0.880 5.320 ;
        RECT -9.010 4.950 -2.830 5.050 ;
        RECT -8.970 4.945 -2.830 4.950 ;
        RECT -11.730 4.915 -11.450 4.945 ;
        RECT -8.970 4.690 -8.170 4.945 ;
        RECT -6.700 4.885 -6.440 4.945 ;
        RECT -12.490 3.845 -5.130 4.110 ;
        RECT -15.585 3.690 -5.130 3.845 ;
        RECT -17.645 1.810 -17.325 2.070 ;
        RECT -17.565 -6.485 -17.410 1.810 ;
        RECT -15.585 0.940 -15.430 3.690 ;
        RECT -12.490 3.630 -5.130 3.690 ;
        RECT -11.665 3.155 -11.510 3.630 ;
        RECT -11.720 2.835 -11.460 3.155 ;
        RECT -3.310 2.440 -2.830 4.945 ;
        RECT -1.820 4.990 -0.880 5.290 ;
        RECT -1.820 3.670 -1.520 4.990 ;
        RECT -1.180 4.960 -0.880 4.990 ;
        RECT -1.840 3.210 -1.360 3.670 ;
        RECT 0.880 3.210 1.360 3.670 ;
        RECT -13.210 0.940 -12.910 2.125 ;
        RECT -5.000 1.960 -2.830 2.440 ;
        RECT -8.400 0.940 -8.100 1.310 ;
        RECT -15.590 0.785 -15.420 0.940 ;
        RECT -13.980 0.855 -6.620 0.940 ;
        RECT -15.585 -2.105 -15.430 0.785 ;
        RECT -14.755 0.565 -6.620 0.855 ;
        RECT -13.980 0.460 -6.620 0.565 ;
        RECT -13.210 0.370 -12.910 0.460 ;
        RECT -5.960 0.040 -5.420 0.520 ;
        RECT -10.370 -0.465 -9.830 -0.435 ;
        RECT -12.820 -0.725 -12.540 -0.695 ;
        RECT -14.760 -0.945 -12.090 -0.725 ;
        RECT -10.630 -0.945 -9.700 -0.465 ;
        RECT -5.855 -0.485 -5.520 0.040 ;
        RECT -5.000 -0.485 -4.520 1.960 ;
        RECT -3.160 0.850 0.980 1.000 ;
        RECT 1.205 0.850 1.360 3.210 ;
        RECT 1.970 0.850 2.125 6.675 ;
        RECT 3.075 3.400 3.335 3.485 ;
        RECT 6.590 3.400 7.070 3.670 ;
        RECT 3.075 3.245 7.070 3.400 ;
        RECT 3.075 3.165 3.335 3.245 ;
        RECT 6.590 3.210 7.070 3.245 ;
        RECT 9.310 3.210 9.790 3.670 ;
        RECT -3.160 0.720 3.735 0.850 ;
        RECT 9.635 0.720 9.790 3.210 ;
        RECT -3.160 0.695 11.980 0.720 ;
        RECT -3.160 0.520 0.980 0.695 ;
        RECT 3.580 0.650 11.980 0.695 ;
        RECT 3.580 0.565 22.570 0.650 ;
        RECT 3.580 0.560 3.735 0.565 ;
        RECT 4.620 0.495 22.570 0.565 ;
        RECT 4.620 0.240 11.980 0.495 ;
        RECT 14.830 0.170 20.350 0.495 ;
        RECT 22.110 0.170 22.570 0.495 ;
        RECT -5.860 -0.635 -4.520 -0.485 ;
        RECT -1.840 -0.635 -1.530 -0.605 ;
        RECT -8.170 -0.745 -7.910 -0.715 ;
        RECT -6.850 -0.745 -6.530 -0.715 ;
        RECT -8.470 -0.945 -6.530 -0.745 ;
        RECT -14.760 -1.270 -14.540 -0.945 ;
        RECT -12.820 -0.975 -12.540 -0.945 ;
        RECT -10.370 -0.975 -9.830 -0.945 ;
        RECT -8.170 -0.975 -7.910 -0.945 ;
        RECT -6.850 -0.975 -6.530 -0.945 ;
        RECT -5.860 -0.885 -1.355 -0.635 ;
        RECT 0.545 -0.660 0.925 -0.630 ;
        RECT 0.300 -0.850 3.970 -0.660 ;
        RECT 11.300 -0.825 11.925 -0.765 ;
        RECT 12.780 -0.820 13.345 -0.120 ;
        RECT 12.730 -0.825 13.345 -0.820 ;
        RECT -5.860 -0.890 -4.520 -0.885 ;
        RECT -5.860 -0.925 -4.530 -0.890 ;
        RECT -1.840 -0.915 -1.530 -0.885 ;
        RECT -5.860 -1.050 -5.570 -0.925 ;
        RECT 0.300 -0.980 5.630 -0.850 ;
        RECT 0.545 -1.010 0.925 -0.980 ;
        RECT 3.640 -0.995 5.630 -0.980 ;
        RECT 7.315 -0.995 7.545 -0.965 ;
        RECT -14.780 -1.590 -14.520 -1.270 ;
        RECT -5.870 -1.470 -5.570 -1.050 ;
        RECT 3.640 -1.165 7.815 -0.995 ;
        RECT 3.640 -1.170 5.630 -1.165 ;
        RECT 7.315 -1.195 7.545 -1.165 ;
        RECT 8.755 -1.255 9.365 -0.885 ;
        RECT 11.300 -1.035 14.020 -0.825 ;
        RECT 15.215 -1.035 15.465 -0.975 ;
        RECT 11.300 -1.225 15.465 -1.035 ;
        RECT 8.755 -1.265 9.145 -1.255 ;
        RECT 11.300 -1.390 14.020 -1.225 ;
        RECT 15.215 -1.285 15.465 -1.225 ;
        RECT 19.090 -1.070 19.405 -1.010 ;
        RECT 19.090 -1.325 23.355 -1.070 ;
        RECT 19.090 -1.390 19.405 -1.325 ;
        RECT 11.300 -1.460 11.925 -1.390 ;
        RECT -5.900 -1.770 -5.540 -1.470 ;
        RECT -13.980 -2.105 -6.620 -1.780 ;
        RECT -3.750 -1.955 -3.490 -1.870 ;
        RECT -3.160 -1.955 0.980 -1.720 ;
        RECT -4.355 -2.045 0.980 -1.955 ;
        RECT -4.355 -2.105 3.615 -2.045 ;
        RECT -15.585 -2.255 -4.205 -2.105 ;
        RECT -3.750 -2.190 -3.490 -2.105 ;
        RECT -3.160 -2.200 3.615 -2.105 ;
        RECT -15.585 -2.260 -6.620 -2.255 ;
        RECT -13.595 -3.510 -13.440 -2.260 ;
        RECT 3.460 -2.280 3.615 -2.200 ;
        RECT 4.620 -2.280 11.980 -2.000 ;
        RECT 12.730 -2.010 13.295 -1.390 ;
        RECT 3.460 -2.325 11.980 -2.280 ;
        RECT 13.495 -2.325 13.650 -2.320 ;
        RECT 14.830 -2.325 20.350 -2.070 ;
        RECT 3.460 -2.395 20.350 -2.325 ;
        RECT 22.110 -2.395 22.570 -2.070 ;
        RECT 3.460 -2.435 22.570 -2.395 ;
        RECT 4.620 -2.480 22.570 -2.435 ;
        RECT -12.030 -3.510 -11.550 -3.400 ;
        RECT -13.595 -3.665 -11.550 -3.510 ;
        RECT -12.030 -3.860 -11.550 -3.665 ;
        RECT -9.310 -3.475 -8.830 -3.400 ;
        RECT -8.210 -3.475 -7.890 -3.420 ;
        RECT 5.280 -3.430 5.580 -2.480 ;
        RECT 13.495 -2.510 13.650 -2.480 ;
        RECT 14.830 -2.550 22.570 -2.480 ;
        RECT -9.310 -3.630 -7.890 -3.475 ;
        RECT 12.700 -3.540 13.325 -2.975 ;
        RECT -9.310 -3.860 -8.830 -3.630 ;
        RECT -8.210 -3.680 -7.890 -3.630 ;
        RECT 12.730 -3.765 13.295 -3.540 ;
        RECT 1.270 -4.330 13.295 -3.765 ;
        RECT 20.650 -4.880 20.795 -2.550 ;
        RECT 5.140 -5.090 5.620 -4.890 ;
        RECT 3.175 -5.245 5.620 -5.090 ;
        RECT 3.175 -5.785 3.330 -5.245 ;
        RECT 5.140 -5.350 5.620 -5.245 ;
        RECT 7.860 -5.350 8.340 -4.890 ;
        RECT 20.650 -5.025 25.170 -4.880 ;
        RECT 3.125 -6.105 3.385 -5.785 ;
        RECT 8.185 -5.855 8.340 -5.350 ;
        RECT -19.205 -6.640 -13.055 -6.485 ;
        RECT -19.205 -6.990 -19.050 -6.640 ;
        RECT -19.490 -7.470 -19.030 -6.990 ;
        RECT -13.210 -7.160 -13.055 -6.640 ;
        RECT -13.700 -7.170 -3.035 -7.160 ;
        RECT -1.000 -7.170 -0.700 -6.140 ;
        RECT 8.135 -6.175 8.395 -5.855 ;
        RECT 8.590 -6.565 8.910 -6.520 ;
        RECT 3.675 -6.735 8.910 -6.565 ;
        RECT 3.675 -6.990 3.845 -6.735 ;
        RECT 8.590 -6.780 8.910 -6.735 ;
        RECT 3.675 -7.075 3.855 -6.990 ;
        RECT 2.510 -7.170 2.830 -7.115 ;
        RECT -13.700 -7.315 2.830 -7.170 ;
        RECT -14.730 -7.380 -14.410 -7.330 ;
        RECT -13.700 -7.380 -6.340 -7.315 ;
        RECT -14.730 -7.535 -6.340 -7.380 ;
        RECT -14.730 -7.590 -14.410 -7.535 ;
        RECT -13.700 -7.640 -6.340 -7.535 ;
        RECT -3.270 -7.325 2.830 -7.315 ;
        RECT -3.270 -7.650 0.870 -7.325 ;
        RECT 2.510 -7.375 2.830 -7.325 ;
        RECT -10.060 -8.535 -9.580 -8.260 ;
        RECT -5.800 -8.450 -5.540 -8.130 ;
        RECT -11.675 -8.825 -11.395 -8.765 ;
        RECT -17.300 -9.045 -11.395 -8.825 ;
        RECT -19.490 -10.035 -19.030 -9.710 ;
        RECT -18.670 -10.035 -18.350 -9.980 ;
        RECT -19.490 -10.190 -18.350 -10.035 ;
        RECT -18.670 -10.240 -18.350 -10.190 ;
        RECT -17.300 -16.160 -17.080 -9.045 ;
        RECT -11.675 -9.105 -11.395 -9.045 ;
        RECT -10.090 -9.075 -9.550 -8.535 ;
        RECT -7.880 -8.845 -7.620 -8.815 ;
        RECT -5.770 -8.845 -5.570 -8.450 ;
        RECT -8.060 -9.045 -5.570 -8.845 ;
        RECT -2.690 -8.805 -2.370 -8.800 ;
        RECT -1.950 -8.805 -1.640 -8.775 ;
        RECT 0.435 -8.800 0.815 -8.770 ;
        RECT -7.880 -9.075 -7.620 -9.045 ;
        RECT -2.690 -9.055 -1.075 -8.805 ;
        RECT 0.320 -8.895 2.380 -8.800 ;
        RECT 3.685 -8.895 3.855 -7.075 ;
        RECT 8.110 -7.170 8.430 -6.925 ;
        RECT 4.120 -7.395 4.380 -7.315 ;
        RECT 4.620 -7.325 13.495 -7.170 ;
        RECT 4.620 -7.395 11.980 -7.325 ;
        RECT 4.120 -7.550 11.980 -7.395 ;
        RECT 4.120 -7.635 4.380 -7.550 ;
        RECT 4.620 -7.650 11.980 -7.550 ;
        RECT 13.340 -7.410 13.495 -7.325 ;
        RECT 14.580 -7.340 20.100 -7.300 ;
        RECT 14.580 -7.410 23.050 -7.340 ;
        RECT 13.340 -7.495 23.050 -7.410 ;
        RECT 13.340 -7.565 20.100 -7.495 ;
        RECT 14.580 -7.780 20.100 -7.565 ;
        RECT 22.590 -7.820 23.050 -7.495 ;
        RECT 13.420 -8.360 13.680 -8.040 ;
        RECT 11.300 -8.510 11.925 -8.455 ;
        RECT 8.680 -8.775 8.850 -8.745 ;
        RECT 5.615 -8.885 5.845 -8.855 ;
        RECT -2.690 -9.060 -2.370 -9.055 ;
        RECT -10.060 -9.390 -9.580 -9.075 ;
        RECT -1.950 -9.085 -1.640 -9.055 ;
        RECT 0.320 -9.065 3.855 -8.895 ;
        RECT 4.215 -9.055 6.075 -8.885 ;
        RECT 0.320 -9.120 2.380 -9.065 ;
        RECT 0.435 -9.150 0.815 -9.120 ;
        RECT 3.510 -9.495 3.830 -9.450 ;
        RECT 4.215 -9.495 4.385 -9.055 ;
        RECT 5.615 -9.085 5.845 -9.055 ;
        RECT 8.585 -9.125 9.025 -8.775 ;
        RECT 11.300 -9.005 12.940 -8.510 ;
        RECT 13.465 -9.005 13.635 -8.360 ;
        RECT 18.855 -8.930 19.110 -8.835 ;
        RECT 18.840 -8.960 19.155 -8.930 ;
        RECT 14.940 -9.005 15.170 -8.975 ;
        RECT 18.735 -8.995 20.105 -8.960 ;
        RECT 11.300 -9.075 15.445 -9.005 ;
        RECT 8.585 -9.145 8.925 -9.125 ;
        RECT 11.300 -9.140 11.925 -9.075 ;
        RECT 8.620 -9.220 8.880 -9.145 ;
        RECT 12.375 -9.175 15.445 -9.075 ;
        RECT -14.705 -9.980 -14.445 -9.660 ;
        RECT 3.510 -9.665 4.385 -9.495 ;
        RECT 3.510 -9.710 3.830 -9.665 ;
        RECT -14.655 -12.820 -14.500 -9.980 ;
        RECT -13.700 -10.120 -6.340 -9.880 ;
        RECT -4.025 -10.120 -3.870 -10.115 ;
        RECT -3.270 -10.120 0.870 -9.890 ;
        RECT 4.620 -10.120 11.980 -9.890 ;
        RECT -13.700 -10.215 11.980 -10.120 ;
        RECT -13.700 -10.275 12.165 -10.215 ;
        RECT -13.700 -10.360 -6.340 -10.275 ;
        RECT -12.890 -11.180 -12.590 -10.360 ;
        RECT -5.090 -11.480 -4.610 -10.740 ;
        RECT -5.075 -11.880 -4.665 -11.480 ;
        RECT -5.110 -12.420 -4.630 -11.880 ;
        RECT -5.000 -12.710 -4.800 -12.420 ;
        RECT -14.655 -12.975 -5.450 -12.820 ;
        RECT -5.000 -12.910 -4.350 -12.710 ;
        RECT -12.810 -13.085 -5.450 -12.975 ;
        RECT -12.810 -13.240 -4.975 -13.085 ;
        RECT -12.810 -13.300 -5.450 -13.240 ;
        RECT -5.130 -13.600 -4.975 -13.240 ;
        RECT -5.215 -13.860 -4.895 -13.600 ;
        RECT -9.200 -14.225 -8.660 -14.195 ;
        RECT -11.655 -14.485 -11.375 -14.455 ;
        RECT -14.750 -14.705 -10.860 -14.485 ;
        RECT -9.450 -14.705 -8.510 -14.225 ;
        RECT -6.985 -14.505 -6.725 -14.475 ;
        RECT -4.550 -14.505 -4.350 -12.910 ;
        RECT -7.620 -14.705 -4.350 -14.505 ;
        RECT -11.655 -14.735 -11.375 -14.705 ;
        RECT -9.200 -14.735 -8.660 -14.705 ;
        RECT -6.985 -14.735 -6.725 -14.705 ;
        RECT -12.810 -15.670 -5.450 -15.540 ;
        RECT -4.025 -15.595 -3.870 -10.275 ;
        RECT -3.270 -10.370 0.870 -10.275 ;
        RECT 4.620 -10.370 12.165 -10.275 ;
        RECT 1.165 -10.960 1.425 -10.640 ;
        RECT 1.215 -11.250 1.370 -10.960 ;
        RECT -1.830 -11.710 -1.350 -11.250 ;
        RECT 0.890 -11.710 1.370 -11.250 ;
        RECT 4.780 -11.000 5.080 -10.970 ;
        RECT 5.380 -11.000 5.680 -10.370 ;
        RECT 12.010 -10.775 12.165 -10.370 ;
        RECT 4.780 -11.300 5.680 -11.000 ;
        RECT 11.960 -11.095 12.220 -10.775 ;
        RECT 4.780 -11.330 5.080 -11.300 ;
        RECT 12.375 -11.720 12.940 -9.175 ;
        RECT 14.940 -9.205 15.170 -9.175 ;
        RECT 18.735 -9.215 23.665 -8.995 ;
        RECT 18.840 -9.225 23.665 -9.215 ;
        RECT 18.840 -9.250 19.425 -9.225 ;
        RECT 18.855 -9.415 19.425 -9.250 ;
        RECT 14.580 -10.260 20.100 -10.020 ;
        RECT 21.650 -10.260 21.795 -10.255 ;
        RECT 22.590 -10.260 23.050 -10.060 ;
        RECT 14.580 -10.360 23.050 -10.260 ;
        RECT 14.010 -10.405 23.050 -10.360 ;
        RECT 14.010 -10.500 20.100 -10.405 ;
        RECT 14.010 -10.580 14.770 -10.500 ;
        RECT 14.010 -10.775 14.230 -10.580 ;
        RECT 13.990 -11.095 14.250 -10.775 ;
        RECT 21.650 -11.475 21.795 -10.405 ;
        RECT 22.590 -10.540 23.050 -10.405 ;
        RECT 25.025 -11.475 25.170 -5.025 ;
        RECT 21.650 -11.620 25.170 -11.475 ;
        RECT 8.530 -11.940 12.990 -11.720 ;
        RECT -2.925 -12.745 -1.770 -12.590 ;
        RECT -2.925 -13.575 -2.770 -12.745 ;
        RECT -2.230 -13.070 -1.770 -12.745 ;
        RECT -2.975 -13.895 -2.715 -13.575 ;
        RECT -2.230 -15.595 -1.770 -15.310 ;
        RECT -4.025 -15.670 -1.770 -15.595 ;
        RECT -12.810 -15.790 -1.770 -15.670 ;
        RECT -12.810 -15.825 -2.015 -15.790 ;
        RECT -12.810 -16.020 -5.450 -15.825 ;
        RECT 8.530 -16.160 8.750 -11.940 ;
        RECT 10.590 -12.000 12.940 -11.940 ;
        RECT -17.300 -16.380 8.750 -16.160 ;
      LAYER met2 ;
        RECT -10.210 7.905 -9.950 7.985 ;
        RECT -13.885 7.750 -9.950 7.905 ;
        RECT -14.755 6.540 -14.405 6.830 ;
        RECT -17.615 2.020 -17.355 2.100 ;
        RECT -16.495 2.020 -16.105 2.095 ;
        RECT -17.615 1.865 -16.105 2.020 ;
        RECT -17.615 1.780 -17.355 1.865 ;
        RECT -16.495 1.795 -16.105 1.865 ;
        RECT -14.725 0.535 -14.435 6.540 ;
        RECT -13.885 3.070 -13.730 7.750 ;
        RECT -10.210 7.665 -9.950 7.750 ;
        RECT -1.210 5.280 -0.850 5.290 ;
        RECT -1.215 5.000 -0.845 5.280 ;
        RECT -1.210 4.990 -0.850 5.000 ;
        RECT 3.130 3.455 3.285 3.685 ;
        RECT 3.045 3.195 3.365 3.455 ;
        RECT -11.750 3.070 -11.430 3.125 ;
        RECT -13.885 2.915 -11.430 3.070 ;
        RECT 3.060 3.060 3.360 3.195 ;
        RECT 3.130 3.015 3.285 3.060 ;
        RECT -11.750 2.865 -11.430 2.915 ;
        RECT -13.200 2.095 -12.920 2.130 ;
        RECT -13.240 1.795 -12.880 2.095 ;
        RECT -13.200 1.760 -12.920 1.795 ;
        RECT -10.210 -0.975 -9.730 2.125 ;
        RECT -2.500 1.850 13.345 2.400 ;
        RECT -4.250 1.835 13.345 1.850 ;
        RECT -4.250 1.370 -1.935 1.835 ;
        RECT -8.390 1.280 -8.110 1.315 ;
        RECT -8.430 0.980 -8.070 1.280 ;
        RECT -8.390 0.945 -8.110 0.980 ;
        RECT -5.930 0.945 -5.450 0.970 ;
        RECT -5.950 0.515 -5.430 0.945 ;
        RECT -5.930 0.010 -5.450 0.515 ;
        RECT -4.250 -0.670 -3.770 1.370 ;
        RECT -2.500 1.330 -1.935 1.370 ;
        RECT 12.780 -0.150 13.345 1.835 ;
        RECT -6.600 -0.685 -3.770 -0.670 ;
        RECT -6.820 -1.005 -3.770 -0.685 ;
        RECT 12.750 -0.715 13.375 -0.150 ;
        RECT -6.600 -1.070 -3.770 -1.005 ;
        RECT -4.250 -1.110 -3.770 -1.070 ;
        RECT 8.950 -1.210 9.210 -0.890 ;
        RECT -14.810 -1.560 -14.490 -1.300 ;
        RECT -14.760 -4.600 -14.540 -1.560 ;
        RECT -5.870 -3.090 -5.570 -1.440 ;
        RECT -3.770 -1.900 -3.470 -1.835 ;
        RECT -3.780 -2.160 -3.460 -1.900 ;
        RECT -3.770 -2.225 -3.470 -2.160 ;
        RECT 8.995 -2.685 9.165 -1.210 ;
        RECT 12.700 -1.980 13.325 -1.415 ;
        RECT 8.850 -2.865 9.165 -2.685 ;
        RECT -5.905 -3.370 -5.535 -3.090 ;
        RECT 4.710 -3.100 4.990 -3.065 ;
        RECT -5.870 -3.380 -5.570 -3.370 ;
        RECT -8.180 -3.400 -7.920 -3.390 ;
        RECT 4.270 -3.400 5.610 -3.100 ;
        RECT 8.850 -3.185 9.035 -2.865 ;
        RECT -8.245 -3.700 -7.855 -3.400 ;
        RECT 4.710 -3.435 4.990 -3.400 ;
        RECT 8.850 -3.500 9.040 -3.185 ;
        RECT -8.180 -3.710 -7.920 -3.700 ;
        RECT 1.390 -4.360 1.955 -3.735 ;
        RECT -14.760 -4.820 -3.930 -4.600 ;
        RECT -5.820 -6.065 -5.520 -5.675 ;
        RECT -14.700 -7.620 -14.440 -7.300 ;
        RECT -14.650 -9.690 -14.495 -7.620 ;
        RECT -5.770 -8.160 -5.570 -6.065 ;
        RECT -5.830 -8.420 -5.510 -8.160 ;
        RECT -10.090 -8.660 -9.550 -8.550 ;
        RECT -10.090 -8.805 -4.310 -8.660 ;
        RECT -4.150 -8.805 -3.930 -4.820 ;
        RECT 1.455 -5.695 1.890 -4.360 ;
        RECT 8.865 -5.345 9.040 -3.500 ;
        RECT 12.730 -3.570 13.295 -1.980 ;
        RECT 8.865 -5.515 13.635 -5.345 ;
        RECT -0.970 -6.170 -0.690 -6.135 ;
        RECT -1.390 -6.470 -0.310 -6.170 ;
        RECT -0.970 -6.505 -0.690 -6.470 ;
        RECT 1.465 -7.565 1.875 -5.695 ;
        RECT 3.095 -6.075 3.415 -5.815 ;
        RECT 3.180 -6.410 3.335 -6.075 ;
        RECT 8.105 -6.145 8.425 -5.885 ;
        RECT 3.110 -6.800 3.410 -6.410 ;
        RECT 8.190 -6.895 8.345 -6.145 ;
        RECT 8.620 -6.810 8.880 -6.490 ;
        RECT 2.540 -7.165 2.800 -7.085 ;
        RECT 2.540 -7.320 4.155 -7.165 ;
        RECT 8.140 -7.215 8.400 -6.895 ;
        RECT 2.540 -7.405 2.800 -7.320 ;
        RECT 4.000 -7.345 4.155 -7.320 ;
        RECT 4.000 -7.555 4.410 -7.345 ;
        RECT -2.660 -8.805 -2.400 -8.770 ;
        RECT -10.090 -8.920 -2.400 -8.805 ;
        RECT -10.090 -9.030 -9.550 -8.920 ;
        RECT -5.055 -9.055 -2.400 -8.920 ;
        RECT -5.055 -9.260 -4.805 -9.055 ;
        RECT -2.660 -9.090 -2.400 -9.055 ;
        RECT -14.735 -9.950 -14.415 -9.690 ;
        RECT -18.640 -10.030 -18.380 -9.950 ;
        RECT -16.195 -10.030 -15.805 -9.955 ;
        RECT -18.640 -10.185 -15.805 -10.030 ;
        RECT -18.640 -10.270 -18.380 -10.185 ;
        RECT -16.195 -10.255 -15.805 -10.185 ;
        RECT -5.090 -10.770 -4.610 -9.260 ;
        RECT 1.485 -9.445 1.855 -7.565 ;
        RECT 4.090 -7.605 4.410 -7.555 ;
        RECT 8.665 -8.930 8.835 -6.810 ;
        RECT 13.465 -8.070 13.635 -5.515 ;
        RECT 13.390 -8.330 13.710 -8.070 ;
        RECT 8.590 -9.190 8.910 -8.930 ;
        RECT 3.540 -9.445 3.800 -9.420 ;
        RECT 1.485 -9.735 3.870 -9.445 ;
        RECT 1.485 -9.775 1.855 -9.735 ;
        RECT 3.540 -9.740 3.800 -9.735 ;
        RECT 1.075 -10.720 1.465 -10.645 ;
        RECT -12.970 -10.850 -12.690 -10.815 ;
        RECT -13.300 -11.150 -12.500 -10.850 ;
        RECT -12.970 -11.185 -12.690 -11.150 ;
        RECT -5.120 -11.250 -4.580 -10.770 ;
        RECT 0.945 -10.875 1.595 -10.720 ;
        RECT 11.930 -10.825 12.250 -10.805 ;
        RECT 13.960 -10.825 14.280 -10.805 ;
        RECT 1.075 -10.945 1.465 -10.875 ;
        RECT 3.880 -11.000 4.160 -10.965 ;
        RECT 3.870 -11.300 5.110 -11.000 ;
        RECT 11.930 -11.045 14.280 -10.825 ;
        RECT 11.930 -11.065 12.250 -11.045 ;
        RECT 13.960 -11.065 14.280 -11.045 ;
        RECT 3.880 -11.335 4.160 -11.300 ;
        RECT -9.020 -12.390 -4.600 -11.910 ;
        RECT -9.020 -14.735 -8.540 -12.390 ;
        RECT -5.185 -13.655 -4.925 -13.570 ;
        RECT -3.005 -13.655 -2.685 -13.605 ;
        RECT -5.185 -13.810 -2.685 -13.655 ;
        RECT -5.185 -13.890 -4.925 -13.810 ;
        RECT -3.005 -13.865 -2.685 -13.810 ;
      LAYER met3 ;
        RECT -1.195 4.975 -0.865 5.305 ;
        RECT -16.475 2.095 -16.125 2.120 ;
        RECT -13.225 2.095 -12.895 2.110 ;
        RECT -16.475 1.795 -12.895 2.095 ;
        RECT -16.475 1.770 -16.125 1.795 ;
        RECT -13.225 1.780 -12.895 1.795 ;
        RECT -10.235 2.080 -9.705 2.105 ;
        RECT -10.235 1.600 -5.450 2.080 ;
        RECT -10.235 1.575 -9.705 1.600 ;
        RECT -8.415 1.290 -8.085 1.295 ;
        RECT -8.415 1.280 -8.020 1.290 ;
        RECT -8.830 0.980 -7.670 1.280 ;
        RECT -8.415 0.970 -8.020 0.980 ;
        RECT -8.415 0.965 -8.085 0.970 ;
        RECT -5.930 0.490 -5.450 1.600 ;
        RECT -1.180 1.400 -0.880 4.975 ;
        RECT 3.060 3.430 3.360 3.680 ;
        RECT 3.035 3.080 3.385 3.430 ;
        RECT -3.770 1.100 -0.880 1.400 ;
        RECT -3.770 -1.855 -3.470 1.100 ;
        RECT -3.795 -2.205 -3.445 -1.855 ;
        RECT -3.770 -2.410 -3.470 -2.205 ;
        RECT -5.885 -3.370 -5.555 -3.065 ;
        RECT 3.060 -3.100 3.360 3.080 ;
        RECT 4.685 -3.100 5.015 -3.085 ;
        RECT -8.225 -3.400 -7.875 -3.375 ;
        RECT -7.130 -3.400 -6.750 -3.390 ;
        RECT -5.885 -3.395 -2.740 -3.370 ;
        RECT -8.570 -3.700 -6.750 -3.400 ;
        RECT -8.225 -3.725 -7.875 -3.700 ;
        RECT -7.130 -3.710 -6.750 -3.700 ;
        RECT -5.870 -3.670 -2.740 -3.395 ;
        RECT 3.060 -3.400 5.015 -3.100 ;
        RECT 4.685 -3.415 5.015 -3.400 ;
        RECT -5.870 -4.800 -5.570 -3.670 ;
        RECT -3.040 -4.300 -2.740 -3.670 ;
        RECT -5.870 -5.270 -5.550 -4.800 ;
        RECT -3.020 -5.270 -2.720 -4.770 ;
        RECT -5.870 -5.400 -2.720 -5.270 ;
        RECT -5.850 -5.570 -2.720 -5.400 ;
        RECT -5.850 -5.720 -5.100 -5.570 ;
        RECT -6.160 -6.020 -5.100 -5.720 ;
        RECT -5.845 -6.045 -5.370 -6.020 ;
        RECT -5.670 -6.050 -5.370 -6.045 ;
        RECT -0.995 -6.170 -0.665 -6.155 ;
        RECT -0.995 -6.470 1.430 -6.170 ;
        RECT 3.110 -6.430 3.410 -6.160 ;
        RECT -0.995 -6.485 -0.665 -6.470 ;
        RECT -16.175 -9.955 -15.825 -9.930 ;
        RECT -16.175 -10.255 -15.190 -9.955 ;
        RECT -16.175 -10.280 -15.825 -10.255 ;
        RECT -15.490 -10.850 -15.190 -10.255 ;
        RECT 1.130 -10.620 1.430 -6.470 ;
        RECT 3.085 -6.780 3.435 -6.430 ;
        RECT 1.095 -10.645 1.445 -10.620 ;
        RECT -12.995 -10.850 -12.665 -10.835 ;
        RECT -15.490 -11.150 -12.665 -10.850 ;
        RECT 0.590 -10.945 1.990 -10.645 ;
        RECT 1.095 -10.970 1.445 -10.945 ;
        RECT -12.995 -11.165 -12.665 -11.150 ;
        RECT 3.110 -11.000 3.410 -6.780 ;
        RECT 3.855 -11.000 4.185 -10.985 ;
        RECT 3.110 -11.300 4.185 -11.000 ;
        RECT 3.855 -11.315 4.185 -11.300 ;
      LAYER met4 ;
        RECT -8.360 1.610 -6.050 1.910 ;
        RECT -8.360 1.295 -8.060 1.610 ;
        RECT -8.375 0.965 -8.045 1.295 ;
        RECT -7.105 -3.400 -6.775 -3.385 ;
        RECT -6.350 -3.400 -6.050 1.610 ;
        RECT -7.440 -3.700 -6.050 -3.400 ;
        RECT -7.105 -3.715 -6.775 -3.700 ;
  END
END layout
END LIBRARY

