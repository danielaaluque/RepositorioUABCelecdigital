magic
tech sky130A
magscale 1 2
timestamp 1760680701
<< nwell >>
rect -1630 1224 -1462 2024
rect -1607 -143 -956 178
rect -1277 -531 -956 -143
rect 12 104 180 772
rect 1704 46 1872 772
rect 3787 -201 4546 120
rect -1896 -852 -956 -531
rect -1277 -862 -956 -852
rect -3812 -1763 -2457 -1442
rect -109 -1765 522 -1444
rect 201 -2386 522 -1765
rect 1410 -1534 1578 -940
rect 3737 -1791 4522 -1470
rect -1373 -2895 -404 -2574
<< pwell >>
rect -1893 1523 -1807 1983
rect -2681 1437 -1807 1523
rect -2679 881 -2597 1437
rect -2679 799 -2281 881
rect -210 402 -126 730
rect -884 318 -126 402
rect -2795 -395 -2613 -201
rect -2795 -577 -2177 -395
rect -884 -262 -800 318
rect 577 571 1561 753
rect 577 -245 759 571
rect -884 -346 -272 -262
rect 577 -427 1107 -245
rect 3905 -387 4511 -301
rect -2359 -767 -2177 -577
rect 1167 -1106 1250 -982
rect 617 -1189 1250 -1106
rect -3883 -2003 -2557 -1821
rect 617 -1884 700 -1189
rect 617 -1967 1019 -1884
rect 3761 -2031 4607 -1849
rect -1273 -3135 -363 -2953
<< locali >>
rect 3044 -245 3049 -211
rect 3087 -245 3109 -211
<< viali >>
rect -2340 989 -2296 1033
rect -1770 989 -1674 1085
rect -1334 989 -1294 1029
rect -2558 -189 -2514 -145
rect -2068 -189 -1972 -93
rect -1628 -189 -1588 -149
rect -362 -177 -312 -127
rect 115 -196 179 -132
rect 1469 -233 1503 -199
rect 1804 -233 1838 -199
rect 2266 -280 2379 -165
rect 3049 -245 3087 -207
rect 3824 -266 3875 -214
rect -2329 -1809 -2285 -1765
rect -2012 -1809 -1916 -1713
rect -1570 -1809 -1530 -1769
rect -384 -1811 -334 -1761
rect 93 -1824 157 -1760
rect 1129 -1811 1163 -1777
rect 1736 -1811 1770 -1777
rect 2266 -1816 2379 -1703
rect 2994 -1835 3028 -1801
rect 3774 -1844 3825 -1792
rect -2325 -2941 -2281 -2897
rect -1834 -2941 -1738 -2845
rect -1391 -2941 -1351 -2901
<< metal1 >>
rect -2032 1591 -2001 1938
rect -2048 1539 -2042 1591
rect -1990 1539 -1984 1591
rect -2945 1366 -2887 1372
rect -2887 1308 -2377 1366
rect -1423 1339 -1392 1965
rect -1105 1335 425 1366
rect -2945 1302 -2887 1308
rect -1804 1086 -1634 1106
rect -1804 1085 -566 1086
rect -2346 1033 -2290 1039
rect -2636 989 -2340 1033
rect -2296 989 -2212 1033
rect -1804 1010 -1770 1085
rect -1802 990 -1770 1010
rect -1794 989 -1770 990
rect -1674 1029 -566 1085
rect -236 1058 -176 1064
rect -1674 989 -1334 1029
rect -1294 989 -566 1029
rect -2346 983 -2290 989
rect -1794 938 -1634 989
rect -1340 977 -1288 989
rect -3117 738 -2373 769
rect -3117 188 -3086 738
rect -2333 631 -2302 749
rect -2344 625 -2292 631
rect -2344 567 -2292 573
rect -662 488 -566 989
rect -364 998 -236 1058
rect -364 716 -304 998
rect -236 992 -176 998
rect -1000 392 -566 488
rect -1680 256 -1620 262
rect -3118 157 -3084 188
rect -3117 -421 -3086 157
rect -2951 113 -2945 171
rect -2887 113 -2563 171
rect -1680 138 -1620 196
rect -1192 8 -1186 104
rect -1090 8 -1084 104
rect -2074 -93 -1966 -87
rect -2564 -145 -2508 -139
rect -2952 -189 -2558 -145
rect -2514 -189 -2418 -145
rect -2126 -189 -2068 -93
rect -1946 -189 -1940 -93
rect -1171 -97 -1104 8
rect -1000 -97 -904 392
rect 241 170 272 685
rect 394 170 425 1335
rect 615 691 667 697
rect 667 649 1349 680
rect 615 633 667 639
rect 67 144 747 170
rect 67 139 955 144
rect 716 113 955 139
rect 716 112 747 113
rect 1927 89 1958 699
rect 2357 99 3000 130
rect 4053 99 4453 130
rect -1172 -127 -904 -97
rect 2556 -30 2669 -24
rect -368 -127 -306 -121
rect -1634 -149 -1582 -143
rect -1370 -149 -1364 -143
rect -1694 -189 -1628 -149
rect -1588 -189 -1364 -149
rect -2952 -254 -2908 -189
rect -2564 -195 -2508 -189
rect -2074 -195 -1966 -189
rect -1634 -195 -1582 -189
rect -1370 -195 -1364 -189
rect -1312 -195 -1306 -143
rect -1172 -177 -362 -127
rect -312 -177 -271 -127
rect 109 -132 185 -126
rect -1172 -178 -904 -177
rect -1172 -185 -906 -178
rect -368 -183 -306 -177
rect -1172 -210 -1114 -185
rect 60 -196 115 -132
rect 179 -170 794 -132
rect 2260 -165 2385 -153
rect 2556 -164 2669 -143
rect 2546 -165 2669 -164
rect 179 -196 1126 -170
rect 1751 -184 1873 -177
rect 109 -202 185 -196
rect 728 -199 1126 -196
rect 1463 -199 1509 -193
rect -2956 -260 -2904 -254
rect -1174 -294 -1114 -210
rect 728 -233 1469 -199
rect 1503 -233 1563 -199
rect 728 -234 1126 -233
rect 1463 -239 1509 -233
rect 1751 -236 1790 -184
rect 1842 -236 1873 -184
rect 1751 -251 1873 -236
rect 1751 -253 1829 -251
rect 2260 -280 2266 -165
rect 2379 -207 2804 -165
rect 3043 -207 3093 -195
rect 2379 -245 3049 -207
rect 3087 -245 3093 -207
rect 2379 -278 2804 -245
rect 3043 -257 3093 -245
rect 3818 -214 3881 -202
rect 3818 -266 3824 -214
rect 3875 -265 4671 -214
rect 3875 -266 3881 -265
rect 3818 -278 3881 -266
rect 2379 -280 2385 -278
rect 2260 -292 2385 -280
rect 2546 -283 2659 -278
rect -2956 -318 -2904 -312
rect -1180 -354 -1174 -294
rect -1114 -354 -1108 -294
rect -750 -380 -698 -374
rect -871 -421 -750 -391
rect -3117 -452 -2749 -421
rect -3821 -659 -3815 -601
rect -3757 -659 -3751 -601
rect -3815 -1297 -3757 -659
rect -2719 -702 -2688 -425
rect -1360 -451 -841 -421
rect -698 -421 -561 -391
rect 2546 -402 2659 -396
rect -750 -438 -698 -432
rect 165 -440 723 -409
rect 692 -456 723 -440
rect 692 -487 991 -456
rect 1056 -620 1116 -444
rect 2699 -465 2730 -464
rect 2362 -496 3015 -465
rect 2699 -502 2730 -496
rect 4017 -510 4453 -479
rect -1642 -695 -1636 -684
rect -3277 -733 -2374 -702
rect -1796 -726 -1636 -695
rect -3277 -1069 -3246 -733
rect -1642 -736 -1636 -726
rect -1584 -736 -1578 -684
rect 1056 -686 1116 -680
rect 2540 -708 2546 -595
rect 2659 -708 2665 -595
rect 2546 -753 2659 -708
rect 254 -866 278 -753
rect 391 -866 2659 -753
rect 635 -1049 1059 -1018
rect -3287 -1075 -3235 -1069
rect -3287 -1133 -3235 -1127
rect 635 -1157 666 -1049
rect 625 -1163 677 -1157
rect 1637 -1171 1668 -1011
rect 625 -1221 677 -1215
rect 1627 -1177 1679 -1171
rect -200 -1234 -140 -1228
rect 1627 -1235 1679 -1229
rect -3841 -1328 -2611 -1297
rect -3841 -1331 -3757 -1328
rect -3841 -1428 -3810 -1331
rect -2642 -1459 -2611 -1328
rect -1349 -1463 -607 -1432
rect -200 -1458 -140 -1294
rect 1718 -1313 1724 -1304
rect 735 -1347 1724 -1313
rect 735 -1398 769 -1347
rect 1718 -1356 1724 -1347
rect 1776 -1356 1782 -1304
rect 735 -1415 771 -1398
rect 502 -1434 508 -1423
rect 140 -1465 508 -1434
rect -2946 -1518 -2940 -1466
rect -2888 -1476 -2882 -1466
rect 502 -1475 508 -1465
rect 560 -1475 566 -1423
rect -2888 -1507 -2681 -1476
rect -2888 -1518 -2882 -1507
rect -1160 -1632 -1108 -1626
rect -2012 -1707 -1916 -1652
rect -1160 -1690 -1108 -1684
rect -2018 -1710 -1910 -1707
rect -2335 -1765 -2279 -1753
rect -3460 -1809 -2329 -1765
rect -2285 -1809 -2279 -1765
rect -3734 -2007 -3728 -1996
rect -3837 -2038 -3728 -2007
rect -3734 -2048 -3728 -2038
rect -3676 -2048 -3670 -1996
rect -3460 -3232 -3416 -1809
rect -2335 -1821 -2279 -1809
rect -2018 -1809 -2012 -1710
rect -1916 -1809 -1910 -1710
rect -1576 -1769 -1524 -1763
rect -1154 -1769 -1114 -1690
rect -1612 -1809 -1570 -1769
rect -1530 -1809 -1114 -1769
rect -2018 -1815 -1910 -1809
rect -1576 -1815 -1524 -1809
rect -538 -1812 -532 -1760
rect -480 -1761 -474 -1760
rect -390 -1761 -328 -1755
rect 87 -1760 163 -1754
rect -480 -1811 -384 -1761
rect -334 -1811 -215 -1761
rect -480 -1812 -474 -1811
rect -2012 -1878 -1916 -1815
rect -390 -1817 -328 -1811
rect 64 -1824 93 -1760
rect 157 -1779 476 -1760
rect 737 -1779 771 -1415
rect 1622 -1437 1628 -1385
rect 1680 -1437 1686 -1385
rect 824 -1469 876 -1463
rect 876 -1510 977 -1479
rect 1639 -1485 1670 -1437
rect 2360 -1465 2699 -1434
rect 2668 -1482 2699 -1465
rect 2668 -1513 2981 -1482
rect 3983 -1499 4565 -1468
rect 824 -1527 876 -1521
rect 2684 -1614 2736 -1608
rect 2684 -1672 2736 -1666
rect 2260 -1702 2385 -1691
rect 2260 -1703 2588 -1702
rect 1736 -1755 1770 -1749
rect 1123 -1777 1169 -1771
rect 1717 -1777 1805 -1755
rect 157 -1813 771 -1779
rect 843 -1811 1129 -1777
rect 1163 -1811 1215 -1777
rect 1717 -1786 1736 -1777
rect 1770 -1786 1805 -1777
rect 157 -1824 476 -1813
rect 87 -1830 163 -1824
rect -2941 -1938 -2889 -1932
rect 702 -1942 708 -1890
rect 760 -1899 766 -1890
rect 843 -1899 877 -1811
rect 1123 -1817 1169 -1811
rect 1717 -1829 1724 -1786
rect 1776 -1825 1805 -1786
rect 2260 -1816 2266 -1703
rect 2379 -1801 2588 -1703
rect 2693 -1801 2727 -1672
rect 3771 -1786 3822 -1767
rect 3768 -1792 3831 -1786
rect 2988 -1801 3034 -1795
rect 2379 -1815 2994 -1801
rect 2379 -1816 2385 -1815
rect 1776 -1829 1785 -1825
rect 2260 -1828 2385 -1816
rect 1724 -1844 1776 -1838
rect 2475 -1835 2994 -1815
rect 3028 -1835 3089 -1801
rect 760 -1933 877 -1899
rect 760 -1942 766 -1933
rect -2941 -1996 -2889 -1990
rect -2931 -2564 -2900 -1996
rect -805 -2024 -774 -2023
rect -2578 -2170 -2518 -2044
rect -1421 -2055 2046 -2024
rect -2578 -2236 -2518 -2230
rect -1018 -2154 -922 -2148
rect -1018 -2296 -922 -2250
rect -1015 -2376 -933 -2296
rect -1022 -2382 -926 -2376
rect -1022 -2484 -926 -2478
rect -1000 -2542 -960 -2484
rect -2931 -2595 -2531 -2564
rect -1000 -2582 -870 -2542
rect -1125 -2648 -995 -2617
rect -1026 -2720 -995 -2648
rect -1043 -2772 -1037 -2720
rect -985 -2772 -979 -2720
rect -1840 -2845 -1732 -2839
rect -2331 -2897 -2275 -2891
rect -2950 -2941 -2325 -2897
rect -2281 -2941 -2172 -2897
rect -1890 -2941 -1834 -2845
rect -1708 -2941 -1702 -2845
rect -1397 -2901 -1345 -2895
rect -910 -2901 -870 -2582
rect -1524 -2941 -1391 -2901
rect -1351 -2941 -870 -2901
rect -2331 -2947 -2275 -2941
rect -1840 -2947 -1732 -2941
rect -1397 -2947 -1345 -2941
rect -805 -3119 -774 -2055
rect 233 -2134 285 -2128
rect 233 -2192 285 -2186
rect 243 -2281 274 -2192
rect 956 -2200 1016 -2194
rect 1076 -2200 1136 -2055
rect 2362 -2074 2433 -2043
rect 2402 -2155 2433 -2074
rect 1016 -2260 1136 -2200
rect 2392 -2161 2444 -2155
rect 2392 -2219 2444 -2213
rect 956 -2266 1016 -2260
rect 2475 -2344 2588 -1835
rect 2988 -1841 3034 -1835
rect 3747 -1843 3774 -1792
rect 3768 -1844 3774 -1843
rect 3825 -1799 4021 -1792
rect 3825 -1844 4733 -1799
rect 3768 -1845 4733 -1844
rect 3768 -1850 3885 -1845
rect 3771 -1883 3885 -1850
rect 2802 -2116 2954 -2072
rect 3928 -2081 4547 -2052
rect 2802 -2155 2846 -2116
rect 2798 -2161 2850 -2155
rect 2798 -2219 2850 -2213
rect 1706 -2388 2598 -2344
rect -585 -2549 -393 -2518
rect -585 -2715 -554 -2549
rect -595 -2721 -543 -2715
rect -595 -2779 -543 -2773
rect -805 -3134 -403 -3119
rect -1309 -3165 -403 -3134
rect 1706 -3232 1750 -2388
rect 2118 -2400 2588 -2388
rect -3460 -3276 1750 -3232
<< via1 >>
rect -2042 1539 -1990 1591
rect -2945 1308 -2887 1366
rect -2344 573 -2292 625
rect -236 998 -176 1058
rect -1680 196 -1620 256
rect -2945 113 -2887 171
rect -1186 8 -1090 104
rect -2042 -189 -1972 -93
rect -1972 -189 -1946 -93
rect 615 639 667 691
rect -1364 -195 -1312 -143
rect 2556 -143 2669 -30
rect -2956 -312 -2904 -260
rect 1790 -199 1842 -184
rect 1790 -233 1804 -199
rect 1804 -233 1838 -199
rect 1838 -233 1842 -199
rect 1790 -236 1842 -233
rect -1174 -354 -1114 -294
rect -3815 -659 -3757 -601
rect -750 -432 -698 -380
rect 2546 -396 2659 -283
rect 1056 -680 1116 -620
rect -1636 -736 -1584 -684
rect 2546 -708 2659 -595
rect 278 -866 391 -753
rect -3287 -1127 -3235 -1075
rect 625 -1215 677 -1163
rect -200 -1294 -140 -1234
rect 1627 -1229 1679 -1177
rect 1724 -1356 1776 -1304
rect -2940 -1518 -2888 -1466
rect 508 -1475 560 -1423
rect -1160 -1684 -1108 -1632
rect -3728 -2048 -3676 -1996
rect -2012 -1713 -1916 -1710
rect -2012 -1806 -1916 -1713
rect -532 -1812 -480 -1760
rect 1628 -1437 1680 -1385
rect 824 -1521 876 -1469
rect 2684 -1666 2736 -1614
rect -2941 -1990 -2889 -1938
rect 708 -1942 760 -1890
rect 1724 -1811 1736 -1786
rect 1736 -1811 1770 -1786
rect 1770 -1811 1776 -1786
rect 1724 -1838 1776 -1811
rect -2578 -2230 -2518 -2170
rect -1018 -2250 -922 -2154
rect -1022 -2478 -926 -2382
rect -1037 -2772 -985 -2720
rect -1804 -2941 -1738 -2845
rect -1738 -2941 -1708 -2845
rect 233 -2186 285 -2134
rect 956 -2260 1016 -2200
rect 2392 -2213 2444 -2161
rect 2798 -2213 2850 -2161
rect -595 -2773 -543 -2721
<< metal2 >>
rect -2042 1591 -1990 1597
rect -2777 1550 -2042 1581
rect -2951 1308 -2945 1366
rect -2887 1308 -2881 1366
rect -2945 311 -2887 1308
rect -2777 614 -2746 1550
rect -2042 1533 -1990 1539
rect -242 1056 -236 1058
rect -176 1056 -170 1058
rect -243 1000 -236 1056
rect -176 1000 -169 1056
rect -242 998 -236 1000
rect -176 998 -170 1000
rect 626 691 657 737
rect 609 681 615 691
rect 667 681 673 691
rect 609 639 612 681
rect 672 639 673 681
rect -2350 614 -2344 625
rect -2777 583 -2344 614
rect -2350 573 -2344 583
rect -2292 573 -2286 625
rect 612 612 672 621
rect 626 603 657 612
rect -3455 253 -2887 311
rect -3815 -601 -3757 -595
rect -3455 -601 -3397 253
rect -2945 171 -2887 253
rect -2945 107 -2887 113
rect -2042 416 -1946 425
rect -500 370 2669 480
rect -2042 -93 -1946 320
rect -850 367 2669 370
rect -850 274 -387 367
rect -1678 256 -1622 263
rect -1686 196 -1680 256
rect -1620 196 -1614 256
rect -1678 189 -1622 196
rect -1186 189 -1090 194
rect -1190 104 -1181 189
rect -1095 104 -1086 189
rect -1190 103 -1186 104
rect -1090 103 -1086 104
rect -1186 2 -1090 8
rect -850 -134 -754 274
rect -500 266 -387 274
rect 2556 -30 2669 367
rect -1320 -137 -754 -134
rect -2042 -195 -1946 -189
rect -1364 -143 -754 -137
rect 2550 -143 2556 -30
rect 2669 -143 2675 -30
rect -1312 -195 -754 -143
rect -1364 -201 -754 -195
rect -1320 -214 -754 -201
rect -850 -222 -754 -214
rect 1790 -184 1842 -178
rect 1790 -242 1842 -236
rect -2962 -312 -2956 -260
rect -2904 -312 -2898 -260
rect -1174 -294 -1114 -288
rect -3757 -659 -3397 -601
rect -3815 -665 -3757 -659
rect -2952 -920 -2908 -312
rect -1174 -500 -1114 -354
rect -754 -376 -694 -367
rect -756 -432 -754 -380
rect -694 -432 -692 -380
rect -754 -445 -694 -436
rect -1174 -560 -362 -500
rect -302 -560 -293 -500
rect 1799 -537 1833 -242
rect 2540 -396 2546 -283
rect 2659 -396 2665 -283
rect -1174 -618 -1114 -560
rect 1770 -573 1833 -537
rect -1181 -674 -1172 -618
rect -1116 -674 -1107 -618
rect 942 -620 998 -613
rect 854 -622 1056 -620
rect 854 -678 942 -622
rect 998 -678 1056 -622
rect -1636 -680 -1584 -678
rect 854 -680 1056 -678
rect 1116 -680 1122 -620
rect 1770 -637 1807 -573
rect 2546 -595 2659 -396
rect -1649 -740 -1640 -680
rect -1580 -740 -1571 -680
rect 942 -687 998 -680
rect 1770 -700 1808 -637
rect -1636 -742 -1584 -740
rect 278 -753 391 -747
rect 278 -872 391 -866
rect -379 -920 -370 -912
rect -2952 -964 -370 -920
rect -1214 -1028 -1078 -1026
rect -3293 -1085 -3287 -1075
rect -3582 -1117 -3287 -1085
rect -3728 -1996 -3676 -1990
rect -3582 -2006 -3550 -1117
rect -3293 -1127 -3287 -1117
rect -3235 -1127 -3229 -1075
rect -1214 -1084 -1170 -1028
rect -1114 -1084 -1078 -1028
rect -1214 -1086 -1078 -1084
rect -1166 -1276 -1117 -1086
rect -2940 -1466 -2888 -1460
rect -2940 -1524 -2888 -1518
rect -2930 -1938 -2899 -1524
rect -1166 -1632 -1114 -1276
rect -1166 -1684 -1160 -1632
rect -1108 -1684 -1102 -1632
rect -2018 -1806 -2012 -1710
rect -1916 -1732 -1910 -1710
rect -1916 -1761 -862 -1732
rect -830 -1761 -786 -964
rect -379 -972 -370 -964
rect -310 -972 -301 -912
rect 291 -1139 378 -872
rect 1773 -1069 1808 -700
rect 2546 -714 2659 -708
rect 1773 -1103 2727 -1069
rect -194 -1234 -138 -1227
rect -278 -1294 -200 -1234
rect -140 -1236 -62 -1234
rect -138 -1292 -62 -1236
rect -140 -1294 -62 -1292
rect -194 -1301 -138 -1294
rect 293 -1513 375 -1139
rect 619 -1215 625 -1163
rect 677 -1215 683 -1163
rect 636 -1282 667 -1215
rect 1621 -1229 1627 -1177
rect 1679 -1229 1685 -1177
rect 622 -1291 682 -1282
rect 622 -1360 682 -1351
rect 1638 -1379 1669 -1229
rect 1724 -1304 1776 -1298
rect 1724 -1362 1776 -1356
rect 1628 -1385 1680 -1379
rect 508 -1423 560 -1417
rect 560 -1464 831 -1433
rect 1628 -1443 1680 -1437
rect 508 -1481 560 -1475
rect 800 -1469 831 -1464
rect 800 -1511 824 -1469
rect -532 -1760 -480 -1754
rect -1916 -1784 -532 -1761
rect -1916 -1806 -1910 -1784
rect -1011 -1811 -532 -1784
rect -1011 -1852 -961 -1811
rect -532 -1818 -480 -1812
rect -2947 -1990 -2941 -1938
rect -2889 -1990 -2883 -1938
rect -3239 -2006 -3230 -1991
rect -3676 -2037 -3230 -2006
rect -3582 -2038 -3550 -2037
rect -3728 -2054 -3676 -2048
rect -3239 -2051 -3230 -2037
rect -3170 -2051 -3161 -1991
rect -1018 -2154 -922 -1852
rect 297 -1889 371 -1513
rect 818 -1521 824 -1511
rect 876 -1521 882 -1469
rect 1733 -1786 1767 -1362
rect 2693 -1614 2727 -1103
rect 2678 -1666 2684 -1614
rect 2736 -1666 2742 -1614
rect 1718 -1838 1724 -1786
rect 1776 -1838 1782 -1786
rect 708 -1889 760 -1884
rect 297 -1890 774 -1889
rect 297 -1942 708 -1890
rect 760 -1942 774 -1890
rect 297 -1947 774 -1942
rect 297 -1955 371 -1947
rect 708 -1948 760 -1947
rect 215 -2144 224 -2129
rect 284 -2134 293 -2129
rect -2594 -2170 -2538 -2163
rect -2660 -2172 -2578 -2170
rect -2660 -2228 -2594 -2172
rect -2660 -2230 -2578 -2228
rect -2518 -2230 -2500 -2170
rect -2594 -2237 -2538 -2230
rect -1024 -2250 -1018 -2154
rect -922 -2250 -916 -2154
rect 189 -2175 224 -2144
rect 215 -2189 224 -2175
rect 285 -2144 293 -2134
rect 285 -2175 319 -2144
rect 285 -2186 293 -2175
rect 284 -2189 293 -2186
rect 776 -2200 832 -2193
rect 774 -2202 956 -2200
rect 774 -2258 776 -2202
rect 832 -2258 956 -2202
rect 774 -2260 956 -2258
rect 1016 -2260 1022 -2200
rect 2386 -2213 2392 -2161
rect 2444 -2165 2450 -2161
rect 2792 -2165 2798 -2161
rect 2444 -2209 2798 -2165
rect 2444 -2213 2450 -2209
rect 2792 -2213 2798 -2209
rect 2850 -2213 2856 -2161
rect 776 -2267 832 -2260
rect -1804 -2478 -1022 -2382
rect -926 -2478 -920 -2382
rect -1804 -2845 -1708 -2478
rect -1037 -2720 -985 -2714
rect -601 -2731 -595 -2721
rect -985 -2762 -595 -2731
rect -1037 -2778 -985 -2772
rect -601 -2773 -595 -2762
rect -543 -2773 -537 -2721
rect -1804 -2947 -1708 -2941
<< via2 >>
rect -234 1000 -178 1056
rect 612 639 615 681
rect 615 639 667 681
rect 667 639 672 681
rect 612 621 672 639
rect -2042 320 -1946 416
rect -1678 198 -1622 254
rect -1181 104 -1095 189
rect -1181 103 -1095 104
rect -754 -380 -694 -376
rect -754 -432 -750 -380
rect -750 -432 -698 -380
rect -698 -432 -694 -380
rect -754 -436 -694 -432
rect -362 -560 -302 -500
rect -1172 -674 -1116 -618
rect 942 -678 998 -622
rect -1640 -684 -1580 -680
rect -1640 -736 -1636 -684
rect -1636 -736 -1584 -684
rect -1584 -736 -1580 -684
rect -1640 -740 -1580 -736
rect -1170 -1084 -1114 -1028
rect -370 -972 -310 -912
rect -194 -1292 -140 -1236
rect -140 -1292 -138 -1236
rect 622 -1351 682 -1291
rect -3230 -2051 -3170 -1991
rect 224 -2134 284 -2129
rect -2594 -2228 -2578 -2172
rect -2578 -2228 -2538 -2172
rect 224 -2186 233 -2134
rect 233 -2186 284 -2134
rect 224 -2189 284 -2186
rect 776 -2258 832 -2202
<< metal3 >>
rect -239 1056 -173 1061
rect -239 1000 -234 1056
rect -178 1000 -173 1056
rect -239 995 -173 1000
rect -2047 416 -1941 421
rect -2047 320 -2042 416
rect -1946 320 -1090 416
rect -2047 315 -1941 320
rect -1683 258 -1617 259
rect -1683 256 -1674 258
rect -1766 254 -1674 256
rect -1610 256 -1604 258
rect -1766 198 -1678 254
rect -1766 196 -1674 198
rect -1683 194 -1674 196
rect -1610 196 -1534 256
rect -1610 194 -1604 196
rect -1683 193 -1617 194
rect -1186 189 -1090 320
rect -236 280 -176 995
rect 612 686 672 736
rect 607 681 677 686
rect 607 621 612 681
rect 672 621 677 681
rect 607 616 677 621
rect -1186 103 -1181 189
rect -1095 103 -1090 189
rect -1186 98 -1090 103
rect -754 220 -176 280
rect -754 -371 -694 220
rect -759 -376 -689 -371
rect -759 -436 -754 -376
rect -694 -436 -689 -376
rect -759 -441 -689 -436
rect -754 -482 -694 -441
rect -367 -500 -297 -495
rect -410 -560 -362 -500
rect -302 -560 -234 -500
rect -374 -565 -297 -560
rect -1176 -613 -1116 -586
rect -1177 -618 -1111 -613
rect -1177 -674 -1172 -618
rect -1116 -674 -1111 -618
rect -374 -624 -314 -565
rect 612 -620 672 616
rect 937 -620 1003 -617
rect 612 -622 1003 -620
rect -1645 -680 -1575 -675
rect -1426 -680 -1420 -678
rect -1714 -740 -1640 -680
rect -1580 -740 -1420 -680
rect -1645 -745 -1575 -740
rect -1426 -742 -1420 -740
rect -1356 -742 -1350 -678
rect -1177 -679 -1096 -674
rect -1176 -734 -1096 -679
rect 612 -678 942 -622
rect 998 -678 1003 -622
rect 612 -680 1003 -678
rect 937 -683 1003 -680
rect -1172 -1023 -1112 -734
rect -375 -912 -305 -832
rect -434 -972 -370 -912
rect -310 -972 -256 -912
rect -375 -977 -305 -972
rect -1175 -1028 -1109 -1023
rect -1175 -1084 -1170 -1028
rect -1114 -1084 -1109 -1028
rect -1175 -1089 -1109 -1084
rect -199 -1234 -133 -1231
rect -199 -1236 286 -1234
rect -199 -1292 -194 -1236
rect -138 -1292 286 -1236
rect 622 -1286 682 -1232
rect -199 -1294 286 -1292
rect -199 -1297 -133 -1294
rect -3235 -1991 -3165 -1986
rect -3235 -2051 -3230 -1991
rect -3170 -2051 -3038 -1991
rect -3235 -2056 -3165 -2051
rect -3098 -2170 -3038 -2051
rect 226 -2124 286 -1294
rect 617 -1291 687 -1286
rect 617 -1351 622 -1291
rect 682 -1351 687 -1291
rect 617 -1356 687 -1351
rect 219 -2129 289 -2124
rect -2599 -2170 -2533 -2167
rect -3098 -2172 -2533 -2170
rect -3098 -2228 -2594 -2172
rect -2538 -2228 -2533 -2172
rect 118 -2189 224 -2129
rect 284 -2189 398 -2129
rect 219 -2194 289 -2189
rect -3098 -2230 -2533 -2228
rect -2599 -2233 -2533 -2230
rect 622 -2200 682 -1356
rect 771 -2200 837 -2197
rect 622 -2202 837 -2200
rect 622 -2258 776 -2202
rect 832 -2258 837 -2202
rect 622 -2260 837 -2258
rect 771 -2263 837 -2260
<< via3 >>
rect -1674 254 -1610 258
rect -1674 198 -1622 254
rect -1622 198 -1610 254
rect -1674 194 -1610 198
rect -1420 -742 -1356 -678
<< metal4 >>
rect -1672 322 -1210 382
rect -1672 259 -1612 322
rect -1675 258 -1609 259
rect -1675 194 -1674 258
rect -1610 194 -1609 258
rect -1675 193 -1609 194
rect -1421 -678 -1355 -677
rect -1421 -680 -1420 -678
rect -1488 -740 -1420 -680
rect -1421 -742 -1420 -740
rect -1356 -680 -1355 -678
rect -1270 -680 -1210 322
rect -1356 -740 -1210 -680
rect -1356 -742 -1355 -740
rect -1421 -743 -1355 -742
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0 ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1760154773
transform 1 0 4518 0 1 -2060
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_1
timestamp 1760154773
transform 0 1 1076 -1 0 -978
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_2
timestamp 1760154773
transform 1 0 4422 0 1 -462
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_3
timestamp 1760154773
transform 1 0 -3898 0 1 -1990
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_4
timestamp 1760154773
transform 0 1 -320 -1 0 734
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_5
timestamp 1760154773
transform 1 0 -446 0 1 -3110
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_6
timestamp 1760154773
transform 0 1 -2358 -1 0 -680
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_7
timestamp 1760154773
transform 0 1 -1984 -1 0 1986
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_8
timestamp 1760154773
transform 0 1 1366 -1 0 734
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_9
timestamp 1760154773
transform 0 1 -318 -1 0 -2250
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_8  x1 ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 -2498 0 1 774
box -38 -48 1510 592
use sky130_fd_sc_hd__nand2_8  x2
timestamp 1704896540
transform 1 0 -2796 0 1 -404
box -38 -48 1510 592
use sky130_fd_sc_hd__nand2_8  x3
timestamp 1704896540
transform 1 0 -2740 0 1 -2024
box -38 -48 1510 592
use sky130_fd_sc_hd__nand2_8  x4
timestamp 1704896540
transform 1 0 -2562 0 1 -3156
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_8  x5 ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 -632 0 1 -392
box -38 -48 866 592
use sky130_fd_sc_hd__inv_8  x6
timestamp 1704896540
transform 1 0 -654 0 1 -2026
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_8  x7 ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 924 0 1 -448
box -38 -48 1510 592
use sky130_fd_sc_hd__nor2_8  x8
timestamp 1704896540
transform 1 0 924 0 1 -2026
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_8  x9 ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 2916 0 1 -2052
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  x10
timestamp 1704896540
transform 1 0 2966 0 1 -462
box -38 -48 1142 592
<< labels >>
rlabel metal1 -2636 989 -2340 1033 7 ENABLE
port 1 w
rlabel metal1 -2950 -2941 -2325 -2897 7 ENABLE
port 2 w
rlabel metal1 3875 -265 4671 -214 3 Qn
port 3 e
rlabel metal1 3825 -1845 4733 -1799 3 Q
port 4 e
rlabel metal1 -3117 738 -2373 769 7 VGND
port 6 w
rlabel metal1 -2887 1308 -2377 1366 7 VPWR
port 5 w
<< end >>
