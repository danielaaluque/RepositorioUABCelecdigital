magic
tech sky130A
magscale 1 2
timestamp 1761871299
<< metal1 >>
rect 25276 30988 25282 31048
rect 25342 30988 25348 31048
rect 16846 26832 16898 26838
rect 16846 26774 16898 26780
rect 16847 25328 16897 26774
rect 20576 25194 20756 25200
rect 18966 25014 20576 25194
rect 20576 25008 20756 25014
rect 16822 24656 16828 24752
rect 16924 24656 17200 24752
rect 25282 24066 25342 30988
rect 25794 27420 25800 27480
rect 25860 27420 25866 27480
rect 24195 24020 25342 24066
rect 13558 23316 13564 23457
rect 13705 23434 15675 23457
rect 13705 23338 16702 23434
rect 13705 23316 15675 23338
rect 25800 22668 25860 27420
rect 24204 22628 25860 22668
rect 19000 21680 19806 21860
rect 19986 21680 19992 21860
rect 16797 21527 16803 21579
rect 16855 21574 16861 21579
rect 16855 21531 17024 21574
rect 16855 21527 16861 21531
<< via1 >>
rect 25282 30988 25342 31048
rect 16846 26780 16898 26832
rect 20576 25014 20756 25194
rect 16828 24656 16924 24752
rect 25800 27420 25860 27480
rect 13564 23316 13705 23457
rect 19806 21680 19986 21860
rect 16803 21527 16855 21579
<< metal2 >>
rect 25802 41862 25858 41869
rect 25800 41860 25860 41862
rect 25800 41804 25802 41860
rect 25858 41804 25860 41860
rect 25282 40910 25342 40912
rect 25275 40854 25284 40910
rect 25340 40854 25349 40910
rect 22142 33236 22202 33238
rect 22135 33180 22144 33236
rect 22200 33180 22209 33236
rect 22142 27291 22202 33180
rect 25282 31048 25342 40854
rect 25282 30982 25342 30988
rect 25800 27480 25860 41804
rect 25800 27414 25860 27420
rect 16847 27241 22203 27291
rect 16847 26832 16897 27241
rect 16840 26780 16846 26832
rect 16898 26780 16904 26832
rect 25805 25194 25975 25198
rect 20570 25014 20576 25194
rect 20756 25189 25980 25194
rect 20756 25019 25805 25189
rect 25975 25019 25980 25189
rect 20756 25014 25980 25019
rect 25805 25010 25975 25014
rect 9088 24597 9097 24812
rect 9312 24804 11452 24812
rect 9312 24777 14064 24804
rect 9312 24752 15695 24777
rect 16828 24752 16924 24758
rect 9312 24656 16828 24752
rect 9312 24631 15695 24656
rect 16828 24650 16924 24656
rect 9312 24604 14064 24631
rect 9312 24597 11452 24604
rect 16273 24280 16333 24289
rect 16273 24211 16333 24220
rect 9380 23287 9389 23485
rect 9587 23457 11965 23485
rect 13564 23457 13705 23463
rect 9587 23316 13564 23457
rect 9587 23287 11965 23316
rect 13564 23310 13705 23316
rect 16281 21575 16324 24211
rect 19806 21860 19986 21866
rect 16803 21579 16855 21585
rect 16281 21532 16803 21575
rect 16803 21521 16855 21527
rect 19806 13119 19986 21680
rect 19802 12949 19811 13119
rect 19981 12949 19990 13119
rect 19806 12944 19986 12949
<< via2 >>
rect 25802 41804 25858 41860
rect 25284 40854 25340 40910
rect 22144 33180 22200 33236
rect 25805 25019 25975 25189
rect 9097 24597 9312 24812
rect 16273 24220 16333 24280
rect 9389 23287 9587 23485
rect 19811 12949 19981 13119
<< metal3 >>
rect 23238 44602 23244 44666
rect 23308 44602 23314 44666
rect 21582 44454 21588 44518
rect 21652 44454 21658 44518
rect 22134 44490 22140 44554
rect 22204 44490 22210 44554
rect 21590 31610 21650 44454
rect 22142 33241 22202 44490
rect 22686 44478 22692 44542
rect 22756 44478 22762 44542
rect 22694 40912 22754 44478
rect 23246 41862 23306 44602
rect 25797 41862 25863 41865
rect 23246 41860 25863 41862
rect 23246 41804 25802 41860
rect 25858 41804 25863 41860
rect 23246 41802 25863 41804
rect 25797 41799 25863 41802
rect 25279 40912 25345 40915
rect 22694 40910 25345 40912
rect 22694 40854 25284 40910
rect 25340 40854 25345 40910
rect 22694 40852 25345 40854
rect 25279 40849 25345 40852
rect 22139 33236 22205 33241
rect 22139 33180 22144 33236
rect 22200 33180 22205 33236
rect 22139 33175 22205 33180
rect 16273 31550 21650 31610
rect 9092 24812 9317 24817
rect 245 24597 251 24812
rect 466 24597 9097 24812
rect 9312 24597 9317 24812
rect 9092 24592 9317 24597
rect 16273 24285 16333 31550
rect 25800 25189 28320 25194
rect 25800 25019 25805 25189
rect 25975 25019 28320 25189
rect 25800 25014 28320 25019
rect 16268 24280 16338 24285
rect 16268 24220 16273 24280
rect 16333 24220 16338 24280
rect 16268 24215 16338 24220
rect 2473 23259 2479 23513
rect 2733 23485 6205 23513
rect 9384 23485 9592 23490
rect 2733 23287 9389 23485
rect 9587 23287 9592 23485
rect 2733 23259 6205 23287
rect 9384 23282 9592 23287
rect 19806 13119 19986 13124
rect 19806 12949 19811 13119
rect 19981 12949 19986 13119
rect 19806 10406 19986 12949
rect 19806 10226 26678 10406
rect 26498 767 26678 10226
rect 28140 4016 28320 25014
rect 28140 3836 30542 4016
rect 30362 1023 30542 3836
rect 30357 845 30363 1023
rect 30541 845 30547 1023
rect 30362 844 30542 845
rect 26493 589 26499 767
rect 26677 589 26683 767
rect 26498 588 26678 589
<< via3 >>
rect 23244 44602 23308 44666
rect 21588 44454 21652 44518
rect 22140 44490 22204 44554
rect 22692 44478 22756 44542
rect 251 24597 466 24812
rect 2479 23259 2733 23513
rect 30363 845 30541 1023
rect 26499 589 26677 767
<< metal4 >>
rect 6134 44952 6194 45152
rect 6686 44952 6746 45152
rect 7238 44952 7298 45152
rect 7790 44952 7850 45152
rect 8342 44952 8402 45152
rect 8894 44952 8954 45152
rect 9446 44952 9506 45152
rect 9998 44952 10058 45152
rect 10550 44952 10610 45152
rect 11102 44952 11162 45152
rect 11654 44952 11714 45152
rect 12206 44952 12266 45152
rect 12758 44952 12818 45152
rect 13310 44952 13370 45152
rect 13862 44952 13922 45152
rect 14414 44952 14474 45152
rect 14966 44952 15026 45152
rect 15518 44952 15578 45152
rect 16070 44952 16130 45152
rect 16622 44952 16682 45152
rect 17174 44952 17234 45152
rect 17726 44952 17786 45152
rect 18278 44952 18338 45152
rect 18830 44952 18890 45152
rect 19382 44952 19442 45152
rect 19934 44952 19994 45152
rect 20486 44952 20546 45152
rect 21038 44952 21098 45152
rect 21590 44519 21650 45152
rect 22142 44555 22202 45152
rect 22139 44554 22205 44555
rect 21587 44518 21653 44519
rect 21587 44454 21588 44518
rect 21652 44454 21653 44518
rect 22139 44490 22140 44554
rect 22204 44490 22205 44554
rect 22694 44543 22754 45152
rect 23246 44667 23306 45152
rect 23798 44952 23858 45152
rect 24350 44952 24410 45152
rect 24902 44952 24962 45152
rect 25454 44952 25514 45152
rect 26006 44952 26066 45152
rect 26558 44952 26618 45152
rect 27110 44952 27170 45152
rect 27662 44952 27722 45152
rect 28214 44952 28274 45152
rect 28766 44952 28826 45152
rect 29318 44952 29378 45152
rect 23243 44666 23309 44667
rect 23243 44602 23244 44666
rect 23308 44602 23309 44666
rect 23243 44601 23309 44602
rect 22139 44489 22205 44490
rect 22691 44542 22757 44543
rect 22691 44478 22692 44542
rect 22756 44478 22757 44542
rect 22691 44477 22757 44478
rect 21587 44453 21653 44454
rect 200 24812 600 44152
rect 200 24597 251 24812
rect 466 24597 600 24812
rect 200 1000 600 24597
rect 800 23513 1200 44152
rect 2478 23513 2734 23514
rect 800 23259 2479 23513
rect 2733 23259 2734 23513
rect 800 1000 1200 23259
rect 2478 23258 2734 23259
rect 30362 1023 30542 1024
rect 30362 845 30363 1023
rect 30541 845 30542 1023
rect 26498 767 26678 768
rect 26498 589 26499 767
rect 26677 589 26678 767
rect 3314 0 3494 200
rect 7178 0 7358 200
rect 11042 0 11222 200
rect 14906 0 15086 200
rect 18770 0 18950 200
rect 22634 0 22814 200
rect 26498 0 26678 589
rect 30362 0 30542 845
use alt  alt_0
timestamp 1761870269
transform 1 0 19768 0 1 24406
box -3162 -3138 4491 1400
<< labels >>
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 29318 44952 29378 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 28214 44952 28274 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 30362 0 30542 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26498 0 26678 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22634 0 22814 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18770 0 18950 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 14906 0 15086 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 11042 0 11222 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 7178 0 7358 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 3314 0 3494 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 27662 44952 27722 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 27110 44952 27170 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 26006 44952 26066 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 25454 44952 25514 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 24902 44952 24962 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 23798 44952 23858 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23246 44952 23306 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22694 44952 22754 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21590 44952 21650 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 21038 44952 21098 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 20486 44952 20546 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 19382 44952 19442 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 9998 44952 10058 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 9446 44952 9506 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 8342 44952 8402 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 7790 44952 7850 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 7238 44952 7298 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 6134 44952 6194 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 14414 44952 14474 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 13862 44952 13922 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 12758 44952 12818 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 12206 44952 12266 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 11654 44952 11714 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 10550 44952 10610 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 18830 44952 18890 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 18278 44952 18338 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 17174 44952 17234 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 16622 44952 16682 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 16070 44952 16130 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 14966 44952 15026 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 600 44152 1 FreeSans 400 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 800 1000 1200 44152 1 FreeSans 400 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
